
--------> /opt/siemens/catapult/2024.1_2-1117371/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_wait_pkg_v1 IS

COMPONENT ccs_in_wait_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    rdy    : OUT std_logic;
    ivld   : OUT std_logic;
    dat    : IN  std_logic_vector(width-1 DOWNTO 0);
    irdy   : IN  std_logic;
    vld    : IN  std_logic
   );
END COMPONENT;

END ccs_in_wait_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_wait_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    rdy   : OUT std_logic;
    ivld  : OUT std_logic;
    dat   : IN  std_logic_vector(width-1 DOWNTO 0);
    irdy  : IN  std_logic;
    vld   : IN  std_logic
  );
END ccs_in_wait_v1;

ARCHITECTURE beh OF ccs_in_wait_v1 IS
  constant stall_const : std_logic := '0';
  SIGNAL stall_ctrl : std_logic;
BEGIN
  stall_ctrl <= stall_const;

  idat <= dat;
  rdy  <= irdy and not stall_ctrl;
  ivld <= vld and not stall_ctrl;

END beh;


--------> /opt/siemens/catapult/2024.1_2-1117371/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_out_wait_pkg_v1 IS

COMPONENT ccs_out_wait_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    dat    : OUT std_logic_vector(width-1 DOWNTO 0);
    irdy   : OUT std_logic;
    vld    : OUT std_logic;
    idat   : IN  std_logic_vector(width-1 DOWNTO 0);
    rdy    : IN  std_logic;
    ivld   : IN  std_logic
  );
END COMPONENT;

END ccs_out_wait_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_out_wait_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    dat   : OUT std_logic_vector(width-1 DOWNTO 0);
    irdy  : OUT std_logic;
    vld   : OUT std_logic;
    idat  : IN  std_logic_vector(width-1 DOWNTO 0);
    rdy   : IN  std_logic;
    ivld  : IN  std_logic
  );
END ccs_out_wait_v1;

ARCHITECTURE beh OF ccs_out_wait_v1 IS
  constant stall_const : std_logic := '0';
  SIGNAL stall_ctrl : std_logic;
BEGIN
  stall_ctrl <= stall_const;

  dat  <= idat;
  irdy <= rdy and not stall_ctrl;
  vld  <= ivld and not stall_ctrl;

END beh;


--------> /opt/siemens/catapult/2024.1_2-1117371/Mgc_home/pkgs/hls_pkgs/src/funcs.vhd 

-- a package of attributes that give verification tools a hint about
-- the function being implemented
PACKAGE attributes IS
  ATTRIBUTE CALYPTO_FUNC : string;
  ATTRIBUTE CALYPTO_DATA_ORDER : string;
end attributes;

-----------------------------------------------------------------------
-- Package that declares synthesizable functions needed for RTL output
-----------------------------------------------------------------------

LIBRARY ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

PACKAGE funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

   FUNCTION maximum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION minimum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2 : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
   
-----------------------------------------------------------------
-- logic functions
-----------------------------------------------------------------

   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION or_v (inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- mux functions
-----------------------------------------------------------------

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC_VECTOR;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- latch functions
-----------------------------------------------------------------
   FUNCTION lat_s(dinput: STD_LOGIC       ; clk: STD_LOGIC; doutput: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- tristate functions
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC       ; control: STD_LOGIC) RETURN STD_LOGIC;
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: SIGNED  ) RETURN STD_LOGIC;

   -- RETURN 2 bits (left => lt, right => eq)
   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED;
 
   FUNCTION fabs(arg1: SIGNED  ) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "**" (l, r: UNSIGNED) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "**" (l, r: SIGNED  ) RETURN SIGNED  ;

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-- *_stdar functions use shift functions from std_logic_arith
-----------------------------------------------------------------

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;

   -----------------------------------------------------------------
   -- *_stdar functions use shift functions from std_logic_arith
   -----------------------------------------------------------------
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC;
   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE;
   --FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR ;

   FUNCTION ceil_log2(size : NATURAL) return NATURAL;
   FUNCTION bits(size : NATURAL) return NATURAL;    

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   
END funcs;


--------------------------- B O D Y ----------------------------


PACKAGE BODY funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC IS
     BEGIN IF arg1 THEN RETURN '1'; ELSE RETURN '0'; END IF; END;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
--     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;

   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
     VARIABLE result: STD_LOGIC_VECTOR(0 DOWNTO 0);
   BEGIN
     result := (0 => arg1);
     RETURN result;
   END;

   FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 > arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION minimum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 < arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;

   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := input1'LENGTH;
     ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
     ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     --synopsys translate_off
     FOR i IN len-1 DOWNTO 0 LOOP
       result(i) := resolved(input1a(i) & input2a(i));
     END LOOP;
     --synopsys translate_on
     RETURN result;
   END;

   FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED) RETURN UNSIGNED IS
   BEGIN RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

   FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED) RETURN SIGNED IS
   BEGIN RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

-----------------------------------------------------------------
-- Logic Functions
-----------------------------------------------------------------

   FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;
   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(and_v(inputs, 1)); END;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(or_v(inputs, 1)); END;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(xor_v(inputs, 1)); END;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result AND inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

   FUNCTION or_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     -- this if is added as a quick fix for a bug in catapult evaluating the loop even if inputs'LENGTH==1
     -- see dts0100971279
     IF icnt2 > 1 THEN
       FOR i IN icnt2-1 DOWNTO 1 LOOP
         inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
         result := result OR inputsx(olenM1 DOWNTO 0);
       END LOOP;
     END IF;
     RETURN result;
   END;

   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result XOR inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

-----------------------------------------------------------------
-- Muxes
-----------------------------------------------------------------
   
   FUNCTION mux_sel2_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(1 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 4;
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector( size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "01" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "10" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "11" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel3_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(2 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 8;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "001" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "010" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "011" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN "100" =>
       result := inputs0(5*size-1 DOWNTO 4*size);
     WHEN "101" =>
       result := inputs0(6*size-1 DOWNTO 5*size);
     WHEN "110" =>
       result := inputs0(7*size-1 DOWNTO 6*size);
     WHEN "111" =>
       result := inputs0(8*size-1 DOWNTO 7*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel4_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(3 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 16;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "0000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "0001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "0010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "0011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "0100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "0101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "0110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "0111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "1000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "1001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "1010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "1011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "1100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "1101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "1110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "1111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel5_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(4 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 32;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0 );
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "00001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "00010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "00011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "00100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "00101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "00110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "00111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "01000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "01001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "01010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "01011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "01100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "01101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "01110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "01111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "10000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "10001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "10010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "10011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "10100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "10101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "10110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "10111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "11000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "11001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "11010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "11011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "11100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "11101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "11110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "11111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel6_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(5 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 64;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "000001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "000010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "000011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "000100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "000101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "000110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "000111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "001000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "001001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "001010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "001011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "001100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "001101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "001110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "001111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "010000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "010001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "010010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "010011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "010100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "010101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "010110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "010111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "011000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "011001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "011010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "011011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "011100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "011101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "011110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "011111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN "100000" =>
       result := inputs0( 33*size-1 DOWNTO 32*size);
     WHEN "100001" =>
       result := inputs0( 34*size-1 DOWNTO 33*size);
     WHEN "100010" =>
       result := inputs0( 35*size-1 DOWNTO 34*size);
     WHEN "100011" =>
       result := inputs0( 36*size-1 DOWNTO 35*size);
     WHEN "100100" =>
       result := inputs0( 37*size-1 DOWNTO 36*size);
     WHEN "100101" =>
       result := inputs0( 38*size-1 DOWNTO 37*size);
     WHEN "100110" =>
       result := inputs0( 39*size-1 DOWNTO 38*size);
     WHEN "100111" =>
       result := inputs0( 40*size-1 DOWNTO 39*size);
     WHEN "101000" =>
       result := inputs0( 41*size-1 DOWNTO 40*size);
     WHEN "101001" =>
       result := inputs0( 42*size-1 DOWNTO 41*size);
     WHEN "101010" =>
       result := inputs0( 43*size-1 DOWNTO 42*size);
     WHEN "101011" =>
       result := inputs0( 44*size-1 DOWNTO 43*size);
     WHEN "101100" =>
       result := inputs0( 45*size-1 DOWNTO 44*size);
     WHEN "101101" =>
       result := inputs0( 46*size-1 DOWNTO 45*size);
     WHEN "101110" =>
       result := inputs0( 47*size-1 DOWNTO 46*size);
     WHEN "101111" =>
       result := inputs0( 48*size-1 DOWNTO 47*size);
     WHEN "110000" =>
       result := inputs0( 49*size-1 DOWNTO 48*size);
     WHEN "110001" =>
       result := inputs0( 50*size-1 DOWNTO 49*size);
     WHEN "110010" =>
       result := inputs0( 51*size-1 DOWNTO 50*size);
     WHEN "110011" =>
       result := inputs0( 52*size-1 DOWNTO 51*size);
     WHEN "110100" =>
       result := inputs0( 53*size-1 DOWNTO 52*size);
     WHEN "110101" =>
       result := inputs0( 54*size-1 DOWNTO 53*size);
     WHEN "110110" =>
       result := inputs0( 55*size-1 DOWNTO 54*size);
     WHEN "110111" =>
       result := inputs0( 56*size-1 DOWNTO 55*size);
     WHEN "111000" =>
       result := inputs0( 57*size-1 DOWNTO 56*size);
     WHEN "111001" =>
       result := inputs0( 58*size-1 DOWNTO 57*size);
     WHEN "111010" =>
       result := inputs0( 59*size-1 DOWNTO 58*size);
     WHEN "111011" =>
       result := inputs0( 60*size-1 DOWNTO 59*size);
     WHEN "111100" =>
       result := inputs0( 61*size-1 DOWNTO 60*size);
     WHEN "111101" =>
       result := inputs0( 62*size-1 DOWNTO 61*size);
     WHEN "111110" =>
       result := inputs0( 63*size-1 DOWNTO 62*size);
     WHEN "111111" =>
       result := inputs0( 64*size-1 DOWNTO 63*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS  --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2 SEVERITY FAILURE;
     --synopsys translate_on
       CASE sel IS
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0( size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1  DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0(size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
       RETURN result;
   END;
--   BEGIN RETURN mux_v(inputs, TO_STDLOGICVECTOR(sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     ALIAS    sel0   : STD_LOGIC_VECTOR( sel'LENGTH-1 DOWNTO 0 ) IS sel;

     VARIABLE sellen : INTEGER RANGE 2-sel'LENGTH TO sel'LENGTH;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2**sel'LENGTH;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
     TYPE inputs_array_type is array(natural range <>) of std_logic_vector( olen - 1 DOWNTO 0);
     VARIABLE inputs_array : inputs_array_type( 2**sel'LENGTH - 1 DOWNTO 0);
   BEGIN
     sellen := sel'LENGTH;
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2**sellen SEVERITY FAILURE;
     sellen := 2-sellen;
     --synopsys translate_on
     CASE sellen IS
     WHEN 1 =>
       CASE sel0(0) IS

       WHEN '1' 
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0(  size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1 DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0( size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
     WHEN 2 =>
       result := mux_sel2_v(inputs, not sel);
     WHEN 3 =>
       result := mux_sel3_v(inputs, not sel);
     WHEN 4 =>
       result := mux_sel4_v(inputs, not sel);
     WHEN 5 =>
       result := mux_sel5_v(inputs, not sel);
     WHEN 6 =>
       result := mux_sel6_v(inputs, not sel);
     WHEN others =>
       -- synopsys translate_off
       IF(Is_X(sel0)) THEN
         result := (others => 'X');
       ELSE
       -- synopsys translate_on
         FOR i in 0 to 2**sel'LENGTH - 1 LOOP
           inputs_array(i) := inputs0( ((i + 1) * olen) - 1  DOWNTO i*olen);
         END LOOP;
         result := inputs_array(CONV_INTEGER( (UNSIGNED(NOT sel0)) ));
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
     END CASE;
     RETURN result;
   END;

 
-----------------------------------------------------------------
-- Latches
-----------------------------------------------------------------

   FUNCTION lat_s(dinput: STD_LOGIC; clk: STD_LOGIC; doutput: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN mux_s(STD_LOGIC_VECTOR'(doutput & dinput), clk); END;

   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR ; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR ) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     --synopsys translate_off
     ASSERT dinput'LENGTH = doutput'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN mux_v(doutput & dinput, clk);
   END;

-----------------------------------------------------------------
-- Tri-States
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC; control: STD_LOGIC) RETURN STD_LOGIC IS
--   BEGIN RETURN TO_STDLOGIC(tri_v(TO_STDLOGICVECTOR(dinput), control)); END;
--
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR ; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
--     VARIABLE result: STD_LOGIC_VECTOR(dinput'range);
--   BEGIN
--     CASE control IS
--     WHEN '0' | 'L' =>
--       result := (others => 'Z');
--     WHEN '1' | 'H' =>
--       FOR i IN dinput'range LOOP
--         result(i) := to_UX01(dinput(i));
--       END LOOP;
--     WHEN others =>
--       -- synopsys translate_off
--       result := (others => 'X');
--       -- synopsys translate_on
--     END CASE;
--     RETURN result;
--   END;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;

   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     VARIABLE diff: UNSIGNED(l'LENGTH DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     diff := ('0'&l) - ('0'&r);
     RETURN diff(l'LENGTH);
   END;
   FUNCTION "<"(l, r: SIGNED  ) RETURN STD_LOGIC IS
   BEGIN
     RETURN (UNSIGNED(l) < UNSIGNED(r)) xor (l(l'LEFT) xor r(r'LEFT));
   END;

   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION "<=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">"(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;
   FUNCTION ">=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;

   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN not or_s(l xor r);
   END;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   --some functions to placate spyglass
   FUNCTION mult_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a*b;
   END mult_natural;

   FUNCTION div_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a/b;
   END div_natural;

   FUNCTION mod_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a mod b;
   END mod_natural;

   FUNCTION add_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a+b;
   END add_unsigned;

   FUNCTION sub_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a-b;
   END sub_unsigned;

   FUNCTION sub_int(a,b : INTEGER) RETURN INTEGER IS
   BEGIN
     return a-b;
   END sub_int;

   FUNCTION concat_0(b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return '0' & b;
   END concat_0;

   FUNCTION concat_uns(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a&b;
   END concat_uns;

   FUNCTION concat_vect(a,b : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     return a&b;
   END concat_vect;





   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED IS
     CONSTANT ninps : NATURAL := arg'LENGTH / width;
     ALIAS    arg0  : UNSIGNED(arg'LENGTH-1 DOWNTO 0) IS arg;
     VARIABLE result: UNSIGNED(width-1 DOWNTO 0);
     VARIABLE from  : INTEGER;
     VARIABLE dto   : INTEGER;
   BEGIN
     --synopsys translate_off
     ASSERT arg'LENGTH = width * ninps SEVERITY FAILURE;
     --synopsys translate_on
     result := (OTHERS => '0');
     FOR i IN ninps-1 DOWNTO 0 LOOP
       --result := result + arg0((i+1)*width-1 DOWNTO i*width);
       from := mult_natural((i+1), width)-1; --2.1.6.3
       dto  := mult_natural(i,width); --2.1.6.3
       result := add_unsigned(result , arg0(from DOWNTO dto) );
     END LOOP;
     RETURN result;
   END faccu;

   FUNCTION  fabs (arg1: SIGNED) RETURN UNSIGNED IS
   BEGIN
     CASE arg1(arg1'LEFT) IS
     WHEN '1'
     --synopsys translate_off
          | 'H'
     --synopsys translate_on
       =>
       RETURN UNSIGNED'("0") - UNSIGNED(arg1);
     WHEN '0'
     --synopsys translate_off
          | 'L'
     --synopsys translate_on
       =>
       RETURN UNSIGNED(arg1);
     WHEN others =>
       RETURN resolve_unsigned(UNSIGNED(arg1), UNSIGNED'("0") - UNSIGNED(arg1));
     END CASE;
   END;

   PROCEDURE divmod(l, r: UNSIGNED; rdiv, rmod: OUT UNSIGNED) IS
     CONSTANT llen: INTEGER := l'LENGTH;
     CONSTANT rlen: INTEGER := r'LENGTH;
     CONSTANT llen_plus_rlen: INTEGER := llen + rlen;
     VARIABLE lbuf: UNSIGNED(llen+rlen-1 DOWNTO 0);
     VARIABLE diff: UNSIGNED(rlen DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT rdiv'LENGTH = llen AND rmod'LENGTH = rlen SEVERITY FAILURE;
     --synopsys translate_on
     lbuf := (others => '0');
     lbuf(llen-1 DOWNTO 0) := l;
     FOR i IN rdiv'range LOOP
       diff := sub_unsigned(lbuf(llen_plus_rlen-1 DOWNTO llen-1) ,(concat_0(r)));
       rdiv(i) := not diff(rlen);
       IF diff(rlen) = '0' THEN
         lbuf(llen_plus_rlen-1 DOWNTO llen-1) := diff;
       END IF;
       lbuf(llen_plus_rlen-1 DOWNTO 1) := lbuf(llen_plus_rlen-2 DOWNTO 0);
     END LOOP;
     rmod := lbuf(llen_plus_rlen-1 DOWNTO llen);
   END divmod;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rdiv;
   END "/";

   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rmod;
   END;

   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN l MOD r; END;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rdiv := UNSIGNED'("0") - rdiv;
     END IF;
     RETURN SIGNED(rdiv); -- overflow problem "1000" / "11"
   END "/";

   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
     CONSTANT rnul: UNSIGNED(r'LENGTH-1 DOWNTO 0) := (others => '0');
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     IF rmod /= rnul AND to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rmod := UNSIGNED(r) + rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "MOD";

   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "REM";

   FUNCTION mult_unsigned(l,r : UNSIGNED) return UNSIGNED is
   BEGIN
     return l*r; 
   END mult_unsigned;

   FUNCTION "**" (l, r : UNSIGNED) RETURN UNSIGNED IS
     CONSTANT llen  : NATURAL := l'LENGTH;
     VARIABLE result: UNSIGNED(llen-1 DOWNTO 0);
     VARIABLE fak   : UNSIGNED(llen-1 DOWNTO 0);
   BEGIN
     fak := l;
     result := (others => '0'); result(0) := '1';
     FOR i IN r'reverse_range LOOP
       --was:result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(result & (result*fak)), r(i)));
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR( concat_uns(result , mult_unsigned(result,fak) )), r(i)));

       fak := mult_unsigned(fak , fak);
     END LOOP;
     RETURN result;
   END "**";

   FUNCTION "**" (l, r : SIGNED) RETURN SIGNED IS
     CONSTANT rlen  : NATURAL := r'LENGTH;
     ALIAS    r0    : SIGNED(0 TO r'LENGTH-1) IS r;
     VARIABLE result: SIGNED(l'range);
   BEGIN
     CASE r(r'LEFT) IS
     WHEN '0'
   --synopsys translate_off
          | 'L'
   --synopsys translate_on
     =>
       result := SIGNED(UNSIGNED(l) ** UNSIGNED(r0(1 TO r'LENGTH-1)));
     WHEN '1'
   --synopsys translate_off
          | 'H'
   --synopsys translate_on
     =>
       result := (others => '0');
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END "**";

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-----------------------------------------------------------------

   FUNCTION add_nat(arg1 : NATURAL; arg2 : NATURAL ) RETURN NATURAL IS
   BEGIN
     return (arg1 + arg2);
   END;
   
--   FUNCTION UNSIGNED_2_BIT_VECTOR(arg1 : NATURAL; arg2 : NATURAL ) RETURN BIT_VECTOR IS
--   BEGIN
--     return (arg1 + arg2);
--   END;
   
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(SIGNED(result), arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
        =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
        =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;


   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     --SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: NATURAL range 1 TO len;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => '0');
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         --was:temp(i2+sw) := result(i2);
         temp_idx := add_nat(i2,sw);
         temp(temp_idx) := result(i2);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: sw_range;
     VARIABLE result_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => sbit);
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         -- was: temp(i2) := result(i2+sw);
         result_idx := add_nat(i2,sw);
         temp(i2) := result(result_idx);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;


   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := arg1'LENGTH;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     VARIABLE temp: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     SUBTYPE sw_range IS NATURAL range 0 TO len-1;
     VARIABLE sw: sw_range;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     result := (others=>'0');
     result := arg1;
     sw := sdir MOD len;
     FOR i IN arg2'reverse_range LOOP
       EXIT WHEN sw = 0;
       IF signd2 AND i = arg2'LEFT THEN 
         sw := sub_int(len,sw); 
       END IF;
       -- temp := result(len-sw-1 DOWNTO 0) & result(len-1 DOWNTO len-sw)
       FOR i2 IN len-1 DOWNTO 0 LOOP
         --was: temp((i2+sw) MOD len) := result(i2);
         temp_idx := add_nat(i2,sw) MOD len;
         temp(temp_idx) := result(i2);
       END LOOP;
       result := mux_v(STD_LOGIC_VECTOR(concat_vect(result,temp)), arg2(i));
       sw := mod_natural(mult_natural(sw,2), len);
     END LOOP;
     RETURN result;
   END frot;

   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, -1); END;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, -1); END;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC IS
     CONSTANT len : INTEGER := vec'LENGTH;
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
   BEGIN
     IF index >= len OR index < 0 THEN
       RETURN 'X';
     END IF;
     RETURN vec0(index);
   END;

   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     CONSTANT indexPwidthM1 : INTEGER := index+width-1; --2.1.6.3
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
     CONSTANT xxx : STD_LOGIC_VECTOR(width-1 DOWNTO 0) := (others => 'X');
   BEGIN
     IF index+width > len OR index < 0 THEN
       RETURN xxx;
     END IF;
     RETURN vec0(indexPwidthM1 DOWNTO index);
   END;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     VARIABLE vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     CONSTANT xxx : STD_LOGIC_VECTOR(len-1 DOWNTO 0) := (others => 'X');
   BEGIN
     vec0 := vec;
     IF index >= len OR index < 0 THEN
       RETURN xxx;
     END IF;
     vec0(index) := dinput;
     RETURN vec0;
   END;

   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE IS
     VARIABLE n_b : POSITIVE;
     VARIABLE p_v : NATURAL;
   BEGIN
     p_v := p;
     FOR i IN 1 TO 32 LOOP
       p_v := div_natural(p_v,2);
       n_b := i;
       EXIT WHEN (p_v = 0);
     END LOOP;
     RETURN n_b;
   END;


--   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
--
--     CONSTANT vlen: INTEGER := vec'LENGTH;
--     CONSTANT ilen: INTEGER := dinput'LENGTH;
--     CONSTANT max_shift: INTEGER := vlen-ilen;
--     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
--     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
--     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
--     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
--     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
--     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
--   BEGIN
--     inp := (others => '0');
--     mask := (others => '0');
--
--     IF index > max_shift OR index < 0 THEN
--       RETURN xxx;
--     END IF;
--
--     shift := CONV_UNSIGNED(index, shift'LENGTH);
--     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
--     mask(ilen-1 DOWNTO 0) := ones;
--     inp := fshl(inp, shift, vlen);
--     mask := fshl(mask, shift, vlen);
--     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
--     RETURN vec0;
--   END;

   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR IS

     type enable_matrix is array (0 to enable'LENGTH-1 ) of std_logic_vector(byte_width-1 downto 0);
     CONSTANT vlen: INTEGER := vec'LENGTH;
     CONSTANT ilen: INTEGER := dinput'LENGTH;
     CONSTANT max_shift: INTEGER := vlen-ilen;
     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask2: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE enables: enable_matrix;
     VARIABLE cat_enables: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0 );
     VARIABLE lsbi : INTEGER;
     VARIABLE msbi : INTEGER;

   BEGIN
     cat_enables := (others => '0');
     lsbi := 0;
     msbi := byte_width-1;
     inp := (others => '0');
     mask := (others => '0');

     IF index > max_shift OR index < 0 THEN
       RETURN xxx;
     END IF;

     --initialize enables
     for i in 0 TO (enable'LENGTH-1) loop
       enables(i)  := (others => enable(i));
       cat_enables(msbi downto lsbi) := enables(i) ;
       lsbi := msbi+1;
       msbi := msbi+byte_width;
     end loop;


     shift := CONV_UNSIGNED(index, shift'LENGTH);
     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
     mask(ilen-1 DOWNTO 0) := UNSIGNED((STD_LOGIC_VECTOR(ones) AND cat_enables));
     inp := fshl(inp, shift, vlen);
     mask := fshl(mask, shift, vlen);
     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
     RETURN vec0;
   END;


   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;
   
   FUNCTION bits(size : NATURAL) return NATURAL is
   begin
     return ceil_log2(size);
   END;

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH) xor conv_std_logic_vector(c, s'LENGTH);
     cout := ( (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH)) or (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) or (conv_std_logic_vector(b, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) );
   END PROCEDURE csa;

   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH);
     cout := (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH));
   END PROCEDURE csha;

END funcs;

--------> /opt/siemens/catapult/2024.1_2-1117371/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_comps.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_comps IS
 
FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
FUNCTION ceil_log2(size : NATURAL) return NATURAL;
 

COMPONENT mgc_not
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_and
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nand
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_or
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xnor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_lut
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_switch
  GENERIC (
    widths  : NATURAL;
    ninps  : NATURAL;
    widtha  : NATURAL;
    ninpa  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(widtha*ninpa - 1 DOWNTO 0);
    c: in  std_logic_vector(widths*ninps - 1 DOWNTO 0);
    s: in  std_logic;
    z: out std_logic_vector(widtha       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux
  GENERIC (
    width  :  NATURAL;
    ctrlw  :  NATURAL;
    p2ctrlw : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width*(2**ctrlw) - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw            - 1 DOWNTO 0);
    z: out std_logic_vector(width            - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux1hot
  GENERIC (
    width  : NATURAL;
    ctrlw  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ctrlw - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw       - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_reg_pos
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;  -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL  -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_reg_neg
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;   -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_generic_reg
  GENERIC(
   width: natural := 8;
   ph_clk: integer range 0 to 1 := 1; -- clock polarity, 1=rising_edge
   ph_en: integer range 0 to 1 := 1;
   ph_a_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   ph_s_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   a_rst_used: integer range 0 to 1 := 1;
   s_rst_used: integer range 0 to 1 := 0;
   en_used: integer range 0 to 1 := 1
  );
  PORT(
   d: std_logic_vector(width-1 downto 0);
   clk: in std_logic;
   en: in std_logic;
   a_rst: in std_logic;
   s_rst: in std_logic;
   q: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_equal
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a : in  std_logic_vector(width-1 DOWNTO 0);
    b : in  std_logic_vector(width-1 DOWNTO 0);
    eq: out std_logic;
    ne: out std_logic
  );
END COMPONENT;

COMPONENT mgc_shift_l
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rot
  GENERIC (
    width  : NATURAL;
    width_s: NATURAL;
    signd_s: NATURAL;      -- 0:unsigned 1:signed
    sleft  : NATURAL;      -- 0:right 1:left;
    log2w  : NATURAL := 0; -- LOG2(width)
    l2wp2  : NATURAL := 0  --2**LOG2(width)
  );
  PORT (
    a : in  std_logic_vector(width  -1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width  -1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_ci
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width_a, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width_a, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width_a,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width_a,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_addc
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_msb
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add3
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_c : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_c : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(ifeqsel(width_c,0,width,width_c)-1 DOWNTO 0);
    d: in  std_logic_vector(0 DOWNTO 0);
    e: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_lt
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic
  );
END COMPONENT;

COMPONENT mgc_add_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_sub_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addc_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     c: in std_logic_vector(0 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addsub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    add: in  std_logic;
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_accu
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_abs
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sqr
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_z : NATURAL    -- <= 2 * width_a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_fast
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_pipe
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 
    s_rst_active  : NATURAL; -- 0 to 1 
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic; --spyglass disable SYNTH_5121,W240
    s_rst : in  std_logic; --spyglass disable SYNTH_5121,W240
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL;
    use_const  : NATURAL
  );
  PORT (
    a   : in  std_logic_vector(width_a-1 DOWNTO 0);
    b   : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0); --spyglass disable SYNTH_5121,W240
    c   : in  std_logic_vector(width_c-1 DOWNTO 0);
    d   : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0); --spyglass disable SYNTH_5121,W240
    cst : in  std_logic_vector(width_e-1 DOWNTO 0); --spyglass disable SYNTH_5121,W240
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2   : NATURAL;
    add_d2   : NATURAL;
    use_const : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2     : in  std_logic_vector(width_b2-1 DOWNTO 0);--spyglass disable SYNTH_5121,W240
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2     : in  std_logic_vector(width_d2-1 DOWNTO 0);--spyglass disable SYNTH_5121,W240
    cst   : in  std_logic_vector(width_e-1 DOWNTO 0);--spyglass disable SYNTH_5121,W240
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;--spyglass disable SYNTH_5121,W240
    s_rst : in  std_logic;--spyglass disable SYNTH_5121,W240
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul4add1
  GENERIC (
    gentype : NATURAL;
    width_a1 : NATURAL;
    signd_a1 : NATURAL;
    width_a2 : NATURAL;
    signd_a2 : NATURAL;
    width_b1 : NATURAL;
    signd_b1 : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c1 : NATURAL;
    signd_c1 : NATURAL;
    width_c2 : NATURAL;
    signd_c2 : NATURAL;
    width_d1 : NATURAL;
    signd_d1 : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    add_a : NATURAL;
    add_b : NATURAL;
    add_c : NATURAL;
    use_const : NATURAL
  );
  PORT (
    a1  : in  std_logic_vector(width_a1-1 DOWNTO 0);
    a2  : in  std_logic_vector(width_a2-1 DOWNTO 0);
    b1  : in  std_logic_vector(width_b1-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c1  : in  std_logic_vector(width_c1-1 DOWNTO 0);
    c2  : in  std_logic_vector(width_c2-1 DOWNTO 0);
    d1  : in  std_logic_vector(width_d1-1 DOWNTO 0);--spyglass disable SYNTH_5121,W240
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);--spyglass disable SYNTH_5121,W240
    c  : in  std_logic_vector(width_c-1 DOWNTO 0); --spyglass disable SYNTH_5121,W240
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul4add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a1 : NATURAL;
    signd_a1 : NATURAL;
    width_a2 : NATURAL;
    signd_a2 : NATURAL;
    width_b1 : NATURAL;
    signd_b1 : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c1 : NATURAL;
    signd_c1 : NATURAL;
    width_c2 : NATURAL;
    signd_c2 : NATURAL;
    width_d1 : NATURAL;
    signd_d1 : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_c  : NATURAL;
    signd_c  : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    add_a : NATURAL;
    add_b : NATURAL;
    add_c : NATURAL;
    use_const : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a1  : in  std_logic_vector(width_a1-1 DOWNTO 0);
    a2  : in  std_logic_vector(width_a2-1 DOWNTO 0);
    b1  : in  std_logic_vector(width_b1-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c1  : in  std_logic_vector(width_c1-1 DOWNTO 0);
    c2  : in  std_logic_vector(width_c2-1 DOWNTO 0);
    d1  : in  std_logic_vector(width_d1-1 DOWNTO 0);--spyglass disable SYNTH_5121,W240
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);--spyglass disable SYNTH_5121,W240
    c   : in  std_logic_vector(width_c-1 DOWNTO 0); --spyglass disable SYNTH_5121,W240
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic; --spyglass disable SYNTH_5121,W240
    s_rst : in  std_logic; --spyglass disable SYNTH_5121,W240
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    use_const : NATURAL
  );
  PORT (
    a:   in  std_logic_vector(width_a-1 DOWNTO 0);
    b:   in  std_logic_vector(width_b-1 DOWNTO 0);
    c:   in  std_logic_vector(width_c-1 DOWNTO 0);
    cst: in  std_logic_vector(width_cst-1 DOWNTO 0); --spyglass disable SYNTH_5121,W240
    d:   in  std_logic_vector(width_d-1 DOWNTO 0); --spyglass disable SYNTH_5121,W240
    z:   out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1_pipe
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    use_const : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_cst-1 DOWNTO 0); --spyglass disable SYNTH_5121,W240
    d     : in  std_logic_vector(width_d-1 DOWNTO 0); --spyglass disable SYNTH_5121,W240
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic; --spyglass disable SYNTH_5121,W240
    s_rst : in  std_logic; --spyglass disable SYNTH_5121,W240
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_cplxmul
  GENERIC (
    width_ar : NATURAL;
    signd_ar : NATURAL;
    width_ai : NATURAL;
    signd_ai : NATURAL;
    width_br : NATURAL;
    signd_br : NATURAL;
    width_bi : NATURAL;
    signd_bi : NATURAL;
    width_zr : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    width_zi : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    add_rr   : NATURAL;
    add_ri   : NATURAL;
    add_ir   : NATURAL;
    add_ii   : NATURAL;
    gentype  : NATURAL
  );
  PORT (
    ar  : in  std_logic_vector(width_ar-1 DOWNTO 0);
    ai  : in  std_logic_vector(width_ai-1 DOWNTO 0);
    br  : in  std_logic_vector(width_br-1 DOWNTO 0);
    bi  : in  std_logic_vector(width_bi-1 DOWNTO 0);
    zr  : out std_logic_vector(width_zr-1 DOWNTO 0);
    zi  : out std_logic_vector(width_zi-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_cplxmul_pipe
  GENERIC (
    width_ar : NATURAL;
    signd_ar : NATURAL;
    width_ai : NATURAL;
    signd_ai : NATURAL;
    width_br : NATURAL;
    signd_br : NATURAL;
    width_bi : NATURAL;
    signd_bi : NATURAL;
    width_zr : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    width_zi : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    add_rr   : NATURAL;
    add_ri   : NATURAL;
    add_ir   : NATURAL;
    add_ii   : NATURAL;
    gentype  : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 --spyglass disable SYNTH_5121,W240
    s_rst_active  : NATURAL; -- 0 to 1 --spyglass disable SYNTH_5121,W240
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    ar  : in  std_logic_vector(width_ar-1 DOWNTO 0);
    ai  : in  std_logic_vector(width_ai-1 DOWNTO 0);
    br  : in  std_logic_vector(width_br-1 DOWNTO 0);
    bi  : in  std_logic_vector(width_bi-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    zr  : out std_logic_vector(width_zr-1 DOWNTO 0);
    zi  : out std_logic_vector(width_zi-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mulacc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_d   : NATURAL;
    is_square: NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0); --spyglass disable SYNTH_5121,W240 
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic; --spyglass disable SYNTH_5121,W240 
    s_rst     : in  std_logic; --spyglass disable SYNTH_5121,W240
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2acc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2: NATURAL;
    signd_b2: NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2: NATURAL;
    signd_d2: NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_cxd : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL;
    square_b: NATURAL;
    square_d: NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2        : in  std_logic_vector(width_b2-1 DOWNTO 0);--spyglass disable SYNTH_5121,W240
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2        : in  std_logic_vector(width_d2-1 DOWNTO 0);--spyglass disable SYNTH_5121,W240
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);--spyglass disable SYNTH_5121,W240
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;--spyglass disable SYNTH_5121,W240
    s_rst     : in  std_logic;--spyglass disable SYNTH_5121,W240
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul4acc_pipe
  GENERIC (
    width_a0 : NATURAL;
    signd_a0 : NATURAL;
    width_a1 : NATURAL;
    signd_a1 : NATURAL;
    width_b0 : NATURAL;
    signd_b0 : NATURAL;
    width_b1 : NATURAL;
    signd_b1 : NATURAL;
    width_c0 : NATURAL;
    signd_c0 : NATURAL;
    width_c1 : NATURAL;
    signd_c1 : NATURAL;
    width_d0 : NATURAL;
    signd_d0 : NATURAL;
    width_d1 : NATURAL;
    signd_d1 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_a : NATURAL;
    add_b : NATURAL;
    add_c : NATURAL;
    min_fb_size : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a0         : in  std_logic_vector(width_a0-1 DOWNTO 0);
    a1         : in  std_logic_vector(width_a1-1 DOWNTO 0);
    b0         : in  std_logic_vector(width_b0-1 DOWNTO 0);
    b1         : in  std_logic_vector(width_b1-1 DOWNTO 0);
    c0         : in  std_logic_vector(width_c0-1 DOWNTO 0);
    c1         : in  std_logic_vector(width_c1-1 DOWNTO 0);
    d0         : in  std_logic_vector(width_d0-1 DOWNTO 0); --spyglass disable SYNTH_5121,W240
    d1         : in  std_logic_vector(width_d1-1 DOWNTO 0); --spyglass disable SYNTH_5121,W240
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);   --spyglass disable SYNTH_5121,W240
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic; --spyglass disable SYNTH_5121,W240
    s_rst     : in  std_logic; --spyglass disable SYNTH_5121,W240
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_div
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mod
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rem
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_csa
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     c: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_csha
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_rom
    GENERIC (
      rom_id : natural := 1;
      size : natural := 33;
      width : natural := 32
      );
    PORT (
      data_in : std_logic_vector((size*width)-1 downto 0);
      addr : std_logic_vector(ceil_log2(size)-1 downto 0);
      data_out : out std_logic_vector(width-1 downto 0)
    );
END COMPONENT;

END mgc_comps;

PACKAGE BODY mgc_comps IS
 
   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;
 
END mgc_comps;

--------> /opt/siemens/catapult/2024.1_2-1117371/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_div IS
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END mgc_div;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

USE work.funcs.all;

ARCHITECTURE beh OF mgc_div IS
BEGIN
  z <= std_logic_vector(unsigned(a) / unsigned(b)) WHEN signd = 0 ELSE
       std_logic_vector(  signed(a) /   signed(b));
END beh;

--------> /opt/siemens/catapult/2024.1_2-1117371/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.vhd 
-- Memory Type:            BLOCK
-- Operating Mode:         Simple Dual Port (2-Port)
-- Clock Mode:             Single Clock
-- 
-- RTL Code RW Resolution: RBW
-- Catapult RW Resolution: RBW
-- 
-- HDL Work Library:       Xilinx_RAMS_lib
-- Component Name:         BLOCK_1R1W_RBW
-- Latency = 1:            RAM with no registers on inputs or outputs
--         = 2:            adds embedded register on RAM output
--         = 3:            adds fabric registers to non-clock input RAM pins
--         = 4:            adds fabric register to output (driven by embedded register from latency=2)
-- suppress_sim_read_addr_range_errs:  0 - report errors  1 - suppress errors

LIBRARY ieee;

  USE ieee.std_logic_1164.all;
  USE ieee.numeric_std.all;
PACKAGE BLOCK_1R1W_RBW_pkg IS
  COMPONENT BLOCK_1R1W_RBW IS
  GENERIC (
    addr_width : integer := 8 ;
    data_width : integer := 7 ;
    depth : integer := 256 ;
    latency : integer := 1 ;
    suppress_sim_read_addr_range_errs : integer := 1 
    
  );
  PORT (
    clk : in std_logic ;
    clken : in std_logic ;
    d : in std_logic_vector(data_width-1 downto 0) ;
    q : out std_logic_vector(data_width-1 downto 0) ;
    radr : in std_logic_vector(addr_width-1 downto 0) ;
    re : in std_logic ;
    wadr : in std_logic_vector(addr_width-1 downto 0) ;
    we : in std_logic 
    
  );
  END COMPONENT;
END BLOCK_1R1W_RBW_pkg;
LIBRARY ieee;

  USE ieee.std_logic_1164.all;
  USE ieee.numeric_std.all;
ENTITY BLOCK_1R1W_RBW IS
  GENERIC (
    addr_width : integer := 8 ;
    data_width : integer := 7 ;
    depth : integer := 256 ;
    latency : integer := 1 ;
    suppress_sim_read_addr_range_errs : integer := 1 
    
  );
  PORT (
    clk : in std_logic ;
    clken : in std_logic ;
    d : in std_logic_vector(data_width-1 downto 0) ;
    q : out std_logic_vector(data_width-1 downto 0) ;
    radr : in std_logic_vector(addr_width-1 downto 0) ;
    re : in std_logic ;
    wadr : in std_logic_vector(addr_width-1 downto 0) ;
    we : in std_logic 
    
  );
 END BLOCK_1R1W_RBW;
ARCHITECTURE rtl OF BLOCK_1R1W_RBW IS
  TYPE ram_t IS ARRAY (depth-1 DOWNTO 0) OF std_logic_vector(data_width-1 DOWNTO 0);
  SIGNAL mem : ram_t := (OTHERS => (OTHERS => '0'));
  ATTRIBUTE ram_style: STRING;
  ATTRIBUTE ram_style OF mem : SIGNAL IS "block";
  ATTRIBUTE syn_ramstyle: STRING;
  ATTRIBUTE syn_ramstyle OF mem : SIGNAL IS "block";
  
  SIGNAL ramq : std_logic_vector(data_width-1 downto 0);
  
BEGIN
-- Port Map
-- readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr READ_ENABLE re
-- writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

-- Access memory with non-registered inputs (latency = 1||2)
  IN_PIN :  IF latency < 3 GENERATE
  BEGIN
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
         IF (clken = '1') THEN
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (suppress_sim_read_addr_range_errs < 1 or to_integer(unsigned(radr)) < depth) THEN
          --pragma translate_on
          ramq <= mem(to_integer(unsigned(radr)));
          --pragma translate_off
          END IF;
          --pragma translate_on
          IF (we = '1') THEN
            mem(to_integer(unsigned(wadr))) <= d;
          END IF;
        END IF;
      END IF;
    END PROCESS;
    
  END GENERATE IN_PIN; 

-- Register all non-clock inputs (latency = 3||4)
  IN_REG :  IF latency > 2 GENERATE
    SIGNAL radr_reg : std_logic_vector(addr_width-1 downto 0);
    SIGNAL re_reg : std_logic;
    SIGNAL d_reg : std_logic_vector(data_width-1 downto 0);
    SIGNAL wadr_reg : std_logic_vector(addr_width-1 downto 0);
    SIGNAL we_reg : std_logic;
    
  BEGIN
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
        IF (clken = '1') THEN
          radr_reg <= radr;
          re_reg <= re;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
        IF (clken = '1') THEN
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        END IF;
      END IF;
    END PROCESS;
    
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
         IF (clken = '1') THEN
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (suppress_sim_read_addr_range_errs < 1 or to_integer(unsigned(radr_reg)) < depth) THEN
          --pragma translate_on
          ramq <= mem(to_integer(unsigned(radr_reg)));
          --pragma translate_off
          END IF;
          --pragma translate_on
          IF (we_reg = '1') THEN
            mem(to_integer(unsigned(wadr_reg))) <= d_reg;
          END IF;
        END IF;
      END IF;
    END PROCESS;
    
  END GENERATE IN_REG;

  out_ram : IF latency = 1 GENERATE
  BEGIN
    q <= ramq;
    
  END GENERATE out_ram;

  out_reg1 : IF ((latency = 2) OR (latency = 3)) GENERATE
    SIGNAL tmpq : std_logic_vector(data_width-1 downto 0);
    
  BEGIN
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
        IF (clken = '1') THEN
          tmpq <= ramq;
        END IF;
      END IF;
    END PROCESS;
    
    q <= tmpq;
    
  END GENERATE out_reg1;

  out_reg2 : IF latency = 4 GENERATE
    SIGNAL tmp1q : std_logic_vector(data_width-1 downto 0);
    
    SIGNAL tmp2q : std_logic_vector(data_width-1 downto 0);
    
  BEGIN
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
        IF (clken = '1') THEN
          tmp1q <= ramq;
        END IF;
      END IF;
    END PROCESS;
    
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
        IF (clken = '1') THEN
          tmp2q <= tmp1q;
        END IF;
      END IF;
    END PROCESS;
    
    q <= tmp2q;
    
  END GENERATE out_reg2;


END rtl;

--------> ./rtl_dutmgc_rom_33_32_20_1.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    2024.1_2/1117371 Production Release
--  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
-- 
--  Generated by:   dr655@ecelinux-16.ece.cornell.edu
--  Generated date: Thu Nov 28 23:23:20 2024
-- ----------------------------------------------------------------------

-- 
LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


PACKAGE dutmgc_rom_33_32_20_1_pkg IS 
  COMPONENT dutmgc_rom_33_32_20_1
    PORT (
      addr : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
    );
  END COMPONENT;
END dutmgc_rom_33_32_20_1_pkg;

PACKAGE BODY dutmgc_rom_33_32_20_1_pkg IS
END dutmgc_rom_33_32_20_1_pkg;

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


USE work.dutmgc_rom_33_32_20_1_pkg.all;
LIBRARY std;

USE std.textio.all;
USE ieee.std_logic_textio.all;

ENTITY dutmgc_rom_33_32_20_1 IS
    PORT (
      addr : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
    );
END dutmgc_rom_33_32_20_1;

ARCHITECTURE v1 OF dutmgc_rom_33_32_20_1 IS
  -- Start of SIF_NL_VHDL::nhl_rom_body
  -- Constants for ROM dimensions
  CONSTANT n_width    : INTEGER := 20;
  CONSTANT n_size     : INTEGER := 32;
  CONSTANT n_addr_w   : INTEGER := 5;
  CONSTANT n_inreg    : INTEGER := 0;
  CONSTANT n_outreg   : INTEGER := 0;
  -- Define data types for ROM storage;
  SUBTYPE  word  IS std_logic_vector((n_width)-1 DOWNTO 0);
  TYPE     lookup_table IS ARRAY (0 to n_size-1) of word;

  SIGNAL mem : lookup_table := lookup_table'(
    word'("11110101111110101010"),
    word'("11111101011111000111"),
    word'("00000011110011011111"),
    word'("11111100010011000010"),
    word'("00110011110001011010"),
    word'("11101110100010111101"),
    word'("11101110111100000110"),
    word'("00010111100010110000"),
    word'("00001000000001000100"),
    word'("00000011101100111101"),
    word'("00000111010101100101"),
    word'("00000100111101011001"),
    word'("00000001100000111110"),
    word'("11100001110001110100"),
    word'("11111100011000010101"),
    word'("11110111011000101010"),
    word'("11011000011011010001"),
    word'("10110011011011110001"),
    word'("11111011110000001111"),
    word'("11110101110011110011"),
    word'("00010011000101001101"),
    word'("11010000000001000001"),
    word'("11111010010111000001"),
    word'("11011110110011011101"),
    word'("11111111100011101111"),
    word'("00001010110111101011"),
    word'("11111110010101011110"),
    word'("00000000111010101100"),
    word'("11011111111101000101"),
    word'("00010011100111010101"),
    word'("00111111100001111001"),
    word'("11111000000011110000")
  );
BEGIN

  -- Reading ROM
  PROCESS(addr)
    VARIABLE idx_addr : INTEGER;
  BEGIN
    idx_addr := conv_integer(unsigned(addr(4 DOWNTO 0)));
    data_out <= mem(idx_addr); --spyglass disable W122 // CAT-35158
  END PROCESS;

END v1;



--------> ./rtl_dutmgc_rom_34_64_8_1.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    2024.1_2/1117371 Production Release
--  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
-- 
--  Generated by:   dr655@ecelinux-16.ece.cornell.edu
--  Generated date: Thu Nov 28 23:23:20 2024
-- ----------------------------------------------------------------------

-- 
LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


PACKAGE dutmgc_rom_34_64_8_1_pkg IS 
  COMPONENT dutmgc_rom_34_64_8_1
    PORT (
      addr : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
  END COMPONENT;
END dutmgc_rom_34_64_8_1_pkg;

PACKAGE BODY dutmgc_rom_34_64_8_1_pkg IS
END dutmgc_rom_34_64_8_1_pkg;

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


USE work.dutmgc_rom_34_64_8_1_pkg.all;
LIBRARY std;

USE std.textio.all;
USE ieee.std_logic_textio.all;

ENTITY dutmgc_rom_34_64_8_1 IS
    PORT (
      addr : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END dutmgc_rom_34_64_8_1;

ARCHITECTURE v1 OF dutmgc_rom_34_64_8_1 IS
  -- Start of SIF_NL_VHDL::nhl_rom_body
  -- Constants for ROM dimensions
  CONSTANT n_width    : INTEGER := 8;
  CONSTANT n_size     : INTEGER := 64;
  CONSTANT n_addr_w   : INTEGER := 6;
  CONSTANT n_inreg    : INTEGER := 0;
  CONSTANT n_outreg   : INTEGER := 0;
  -- Define data types for ROM storage;
  SUBTYPE  word  IS std_logic_vector((n_width)-1 DOWNTO 0);
  TYPE     lookup_table IS ARRAY (0 to n_size-1) of word;

  SIGNAL mem : lookup_table := lookup_table'(
    word'("10010010"),
    word'("00100101"),
    word'("10100110"),
    word'("01100001"),
    word'("10100101"),
    word'("00100000"),
    word'("01100001"),
    word'("00000100"),
    word'("01010001"),
    word'("00010100"),
    word'("10100101"),
    word'("01010101"),
    word'("10001000"),
    word'("10010110"),
    word'("10100000"),
    word'("00011010"),
    word'("01001001"),
    word'("10100010"),
    word'("01011001"),
    word'("10101010"),
    word'("10100010"),
    word'("10100110"),
    word'("00100100"),
    word'("10100100"),
    word'("00100110"),
    word'("10100010"),
    word'("01000000"),
    word'("00010100"),
    word'("00101001"),
    word'("10011001"),
    word'("00000010"),
    word'("01100010"),
    word'("10000110"),
    word'("01011010"),
    word'("10000100"),
    word'("01010000"),
    word'("01101010"),
    word'("01011000"),
    word'("01000000"),
    word'("00100001"),
    word'("01101001"),
    word'("01010110"),
    word'("10100110"),
    word'("01000000"),
    word'("01010001"),
    word'("01101001"),
    word'("01100100"),
    word'("00011001"),
    word'("00000001"),
    word'("10010100"),
    word'("01101000"),
    word'("00001001"),
    word'("00010001"),
    word'("00010000"),
    word'("00100100"),
    word'("10000000"),
    word'("00000000"),
    word'("00011010"),
    word'("01010110"),
    word'("00010101"),
    word'("00001000"),
    word'("00001010"),
    word'("00101000"),
    word'("00101010")
  );
BEGIN

  -- Reading ROM
  PROCESS(addr)
    VARIABLE idx_addr : INTEGER;
  BEGIN
    idx_addr := conv_integer(unsigned(addr(5 DOWNTO 0)));
    data_out <= mem(idx_addr); --spyglass disable W122 // CAT-35158
  END PROCESS;

END v1;



--------> ./rtl_dutmgc_rom_35_64_8_1.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    2024.1_2/1117371 Production Release
--  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
-- 
--  Generated by:   dr655@ecelinux-16.ece.cornell.edu
--  Generated date: Thu Nov 28 23:23:20 2024
-- ----------------------------------------------------------------------

-- 
LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


PACKAGE dutmgc_rom_35_64_8_1_pkg IS 
  COMPONENT dutmgc_rom_35_64_8_1
    PORT (
      addr : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
  END COMPONENT;
END dutmgc_rom_35_64_8_1_pkg;

PACKAGE BODY dutmgc_rom_35_64_8_1_pkg IS
END dutmgc_rom_35_64_8_1_pkg;

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


USE work.dutmgc_rom_35_64_8_1_pkg.all;
LIBRARY std;

USE std.textio.all;
USE ieee.std_logic_textio.all;

ENTITY dutmgc_rom_35_64_8_1 IS
    PORT (
      addr : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END dutmgc_rom_35_64_8_1;

ARCHITECTURE v1 OF dutmgc_rom_35_64_8_1 IS
  -- Start of SIF_NL_VHDL::nhl_rom_body
  -- Constants for ROM dimensions
  CONSTANT n_width    : INTEGER := 8;
  CONSTANT n_size     : INTEGER := 64;
  CONSTANT n_addr_w   : INTEGER := 6;
  CONSTANT n_inreg    : INTEGER := 0;
  CONSTANT n_outreg   : INTEGER := 0;
  -- Define data types for ROM storage;
  SUBTYPE  word  IS std_logic_vector((n_width)-1 DOWNTO 0);
  TYPE     lookup_table IS ARRAY (0 to n_size-1) of word;

  SIGNAL mem : lookup_table := lookup_table'(
    word'("10010110"),
    word'("01101001"),
    word'("10101000"),
    word'("10100101"),
    word'("10000110"),
    word'("10100100"),
    word'("10011001"),
    word'("01100110"),
    word'("10100101"),
    word'("01010010"),
    word'("00000010"),
    word'("01010101"),
    word'("00000010"),
    word'("01010110"),
    word'("01000010"),
    word'("10010110"),
    word'("00010110"),
    word'("01010110"),
    word'("00000101"),
    word'("00011010"),
    word'("01101000"),
    word'("01010100"),
    word'("00011010"),
    word'("01010101"),
    word'("10011010"),
    word'("01100101"),
    word'("00000101"),
    word'("01010010"),
    word'("10010001"),
    word'("00010000"),
    word'("01000101"),
    word'("00010101"),
    word'("00011000"),
    word'("01010110"),
    word'("00001001"),
    word'("01000001"),
    word'("01010110"),
    word'("01001010"),
    word'("01101001"),
    word'("10000110"),
    word'("10101010"),
    word'("10000100"),
    word'("10100110"),
    word'("00011000"),
    word'("01011001"),
    word'("00100001"),
    word'("10000100"),
    word'("10011010"),
    word'("10010110"),
    word'("10101010"),
    word'("01001000"),
    word'("00100001"),
    word'("01010001"),
    word'("00101000"),
    word'("01101000"),
    word'("01001001"),
    word'("10000110"),
    word'("01001001"),
    word'("10010110"),
    word'("10100101"),
    word'("10011000"),
    word'("10000110"),
    word'("10100101"),
    word'("01000100")
  );
BEGIN

  -- Reading ROM
  PROCESS(addr)
    VARIABLE idx_addr : INTEGER;
  BEGIN
    idx_addr := conv_integer(unsigned(addr(5 DOWNTO 0)));
    data_out <= mem(idx_addr); --spyglass disable W122 // CAT-35158
  END PROCESS;

END v1;



--------> ./rtl_dutmgc_rom_36_960_15_1.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    2024.1_2/1117371 Production Release
--  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
-- 
--  Generated by:   dr655@ecelinux-16.ece.cornell.edu
--  Generated date: Thu Nov 28 23:23:20 2024
-- ----------------------------------------------------------------------

-- 
LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


PACKAGE dutmgc_rom_36_960_15_1_pkg IS 
  COMPONENT dutmgc_rom_36_960_15_1
    PORT (
      addr : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(14 DOWNTO 0)
    );
  END COMPONENT;
END dutmgc_rom_36_960_15_1_pkg;

PACKAGE BODY dutmgc_rom_36_960_15_1_pkg IS
END dutmgc_rom_36_960_15_1_pkg;

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


USE work.dutmgc_rom_36_960_15_1_pkg.all;
LIBRARY std;

USE std.textio.all;
USE ieee.std_logic_textio.all;

ENTITY dutmgc_rom_36_960_15_1 IS
    PORT (
      addr : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(14 DOWNTO 0)
    );
END dutmgc_rom_36_960_15_1;

ARCHITECTURE v1 OF dutmgc_rom_36_960_15_1 IS
  -- Start of SIF_NL_VHDL::nhl_rom_body
  -- Constants for ROM dimensions
  CONSTANT n_width    : INTEGER := 15;
  CONSTANT n_size     : INTEGER := 960;
  CONSTANT n_addr_w   : INTEGER := 10;
  CONSTANT n_inreg    : INTEGER := 0;
  CONSTANT n_outreg   : INTEGER := 0;
  -- Define data types for ROM storage;
  SUBTYPE  word  IS std_logic_vector((n_width)-1 DOWNTO 0);
  TYPE     lookup_table IS ARRAY (0 to n_size-1) of word;

  SIGNAL mem : lookup_table := lookup_table'(
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("100010100110001"),
    word'("101011011001100"),
    word'("110001101111111"),
    word'("110110001001110"),
    word'("111001001101011"),
    word'("111011010110010"),
    word'("111100110101111"),
    word'("111101110110100"),
    word'("111110100010100"),
    word'("111110111110110"),
    word'("111111010011111"),
    word'("111111100011111"),
    word'("111111101011000"),
    word'("111111110000000"),
    word'("111111110101000"),
    word'("111111111011000"),
    word'("111111111011001"),
    word'("111111111101111"),
    word'("111111111111111"),
    word'("111111111101001"),
    word'("111111111110000"),
    word'("111111111110101"),
    word'("111111111111000"),
    word'("111111111111011"),
    word'("111111111111100"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("100010100110001"),
    word'("101011011001100"),
    word'("110001101111111"),
    word'("110110001001110"),
    word'("111001001101011"),
    word'("111011010110010"),
    word'("111100110101111"),
    word'("111101110110100"),
    word'("111110100010100"),
    word'("111110111110110"),
    word'("111111010011111"),
    word'("111111100011111"),
    word'("111111101011000"),
    word'("111111110000000"),
    word'("111111110101000"),
    word'("111111111011000"),
    word'("111111111011001"),
    word'("111111111101111"),
    word'("111111111111111"),
    word'("111111111101001"),
    word'("111111111110000"),
    word'("111111111110101"),
    word'("111111111111000"),
    word'("111111111111011"),
    word'("111111111111100"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("000000000000000"),
    word'("100101010110111"),
    word'("111010111000101"),
    word'("001101001111100"),
    word'("011011100100001"),
    word'("100110010101000"),
    word'("101110000111001"),
    word'("110011101000001"),
    word'("110111011101001"),
    word'("111010001011001"),
    word'("111011111111001"),
    word'("111101010001110"),
    word'("111110001000101"),
    word'("111110101100110"),
    word'("111111001000101"),
    word'("111111011000000"),
    word'("111111100100001"),
    word'("111111101100101"),
    word'("111111110011111"),
    word'("111111110111101"),
    word'("111111111000110"),
    word'("111111111100011"),
    word'("111111111110110"),
    word'("111111111100011"),
    word'("111111111101100"),
    word'("111111111110010"),
    word'("111111111110111"),
    word'("111111111111001"),
    word'("111111111111011"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("000000000000000"),
    word'("100101010110111"),
    word'("111010111000101"),
    word'("001101001111100"),
    word'("011011100100001"),
    word'("100110010101000"),
    word'("101110000111001"),
    word'("110011101000001"),
    word'("110111011101001"),
    word'("111010001011001"),
    word'("111011111111001"),
    word'("111101010001110"),
    word'("111110001000101"),
    word'("111110101100110"),
    word'("111111001000101"),
    word'("111111011000000"),
    word'("111111100100001"),
    word'("111111101100101"),
    word'("111111110011111"),
    word'("111111110111101"),
    word'("111111111000110"),
    word'("111111111100011"),
    word'("111111111110110"),
    word'("111111111100011"),
    word'("111111111101100"),
    word'("111111111110010"),
    word'("111111111110111"),
    word'("111111111111001"),
    word'("111111111111011"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("000000000000000"),
    word'("000000101001111"),
    word'("001101101010101"),
    word'("100010110110100"),
    word'("111000100010001"),
    word'("001011010110001"),
    word'("011010001100100"),
    word'("100101010011001"),
    word'("101101010110101"),
    word'("110011000111100"),
    word'("110111000101010"),
    word'("111001111011000"),
    word'("111011110100110"),
    word'("111101001010010"),
    word'("111110000010010"),
    word'("111110101001100"),
    word'("111111000111101"),
    word'("111111011000101"),
    word'("111111100101111"),
    word'("111111101111001"),
    word'("111111110010111"),
    word'("111111110110111"),
    word'("111111111000010"),
    word'("111111111100000"),
    word'("111111111110100"),
    word'("111111111100010"),
    word'("111111111101011"),
    word'("111111111110010"),
    word'("111111111110110"),
    word'("111111111111001"),
    word'("111111111111011"),
    word'("111111111111101"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("000000101001111"),
    word'("001101101010101"),
    word'("100010110110100"),
    word'("111000100010001"),
    word'("001011010110001"),
    word'("011010001100100"),
    word'("100101010011001"),
    word'("101101010110101"),
    word'("110011000111100"),
    word'("110111000101010"),
    word'("111001111011000"),
    word'("111011110100110"),
    word'("111101001010010"),
    word'("111110000010010"),
    word'("111110101001100"),
    word'("111111000111101"),
    word'("111111011000101"),
    word'("111111100101111"),
    word'("111111101111001"),
    word'("111111110010111"),
    word'("111111110110111"),
    word'("111111111000010"),
    word'("111111111100000"),
    word'("111111111110100"),
    word'("111111111100010"),
    word'("111111111101011"),
    word'("111111111110010"),
    word'("111111111110110"),
    word'("111111111111001"),
    word'("111111111111011"),
    word'("111111111111101"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("010110001001010"),
    word'("000000110011100"),
    word'("000101011101111"),
    word'("010111110010000"),
    word'("101101111111101"),
    word'("000010011111111"),
    word'("010011010000111"),
    word'("100000001011000"),
    word'("101001101001011"),
    word'("110000011100111"),
    word'("110101010001000"),
    word'("111000101000101"),
    word'("111010111101101"),
    word'("111100100001110"),
    word'("111101101001110"),
    word'("111110011001100"),
    word'("111110111011001"),
    word'("111111010000000"),
    word'("111111011110100"),
    word'("111111101011010"),
    word'("111111110001100"),
    word'("111111110111010"),
    word'("111111111001111"),
    word'("111111111010011"),
    word'("111111111101011"),
    word'("111111111111100"),
    word'("111111111100111"),
    word'("111111111101111"),
    word'("111111111110100"),
    word'("111111111111000"),
    word'("111111111111010"),
    word'("111111111111100"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("010110001001010"),
    word'("000000110011100"),
    word'("000101011101111"),
    word'("010111110010000"),
    word'("101101111111101"),
    word'("000010011111111"),
    word'("010011010000111"),
    word'("100000001011000"),
    word'("101001101001011"),
    word'("110000011100111"),
    word'("110101010001000"),
    word'("111000101000101"),
    word'("111010111101101"),
    word'("111100100001110"),
    word'("111101101001110"),
    word'("111110011001100"),
    word'("111110111011001"),
    word'("111111010000000"),
    word'("111111011110100"),
    word'("111111101011010"),
    word'("111111110001100"),
    word'("111111110111010"),
    word'("111111111001111"),
    word'("111111111010011"),
    word'("111111111101011"),
    word'("111111111111100"),
    word'("111111111100111"),
    word'("111111111101111"),
    word'("111111111110100"),
    word'("111111111111000"),
    word'("111111111111010"),
    word'("111111111111100"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("010010001011110"),
    word'("011100100110101"),
    word'("000010001100001"),
    word'("000011011011100"),
    word'("010100011001011"),
    word'("101010011001011"),
    word'("111111010101111"),
    word'("010000110100011"),
    word'("011110010100110"),
    word'("101000010100101"),
    word'("101111100000100"),
    word'("110100100110010"),
    word'("111000001001101"),
    word'("111010101000100"),
    word'("111100010101011"),
    word'("111101011110001"),
    word'("111110010000010"),
    word'("111110110110010"),
    word'("111111001101110"),
    word'("111111011110010"),
    word'("111111101000100"),
    word'("111111101111101"),
    word'("111111110101111"),
    word'("111111111000111"),
    word'("111111111001110"),
    word'("111111111101000"),
    word'("111111111111001"),
    word'("111111111100110"),
    word'("111111111101110"),
    word'("111111111110011"),
    word'("111111111110111"),
    word'("111111111111010"),
    word'("111111111111100"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("010010001011110"),
    word'("011100100110101"),
    word'("000010001100001"),
    word'("000011011011100"),
    word'("010100011001011"),
    word'("101010011001011"),
    word'("111111010101111"),
    word'("010000110100011"),
    word'("011110010100110"),
    word'("101000010100101"),
    word'("101111100000100"),
    word'("110100100110010"),
    word'("111000001001101"),
    word'("111010101000100"),
    word'("111100010101011"),
    word'("111101011110001"),
    word'("111110010000010"),
    word'("111110110110010"),
    word'("111111001101110"),
    word'("111111011110010"),
    word'("111111101000100"),
    word'("111111101111101"),
    word'("111111110101111"),
    word'("111111111000111"),
    word'("111111111001110"),
    word'("111111111101000"),
    word'("111111111111001"),
    word'("111111111100110"),
    word'("111111111101110"),
    word'("111111111110011"),
    word'("111111111110111"),
    word'("111111111111010"),
    word'("111111111111100"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111101011101101"),
    word'("001111001001100"),
    word'("011010100011101"),
    word'("000001101110001"),
    word'("000100000000010"),
    word'("010101011100000"),
    word'("101011011111000"),
    word'("000000010011111"),
    word'("010001100100101"),
    word'("011110111001101"),
    word'("101000110001001"),
    word'("101111110101001"),
    word'("110100110101110"),
    word'("111000010100001"),
    word'("111010101101010"),
    word'("111100011001111"),
    word'("111101100000010"),
    word'("111110010100101"),
    word'("111110110101000"),
    word'("111111001111101"),
    word'("111111011111101"),
    word'("111111101001011"),
    word'("111111110000001"),
    word'("111111110110010"),
    word'("111111111001010"),
    word'("111111111001111"),
    word'("111111111101001"),
    word'("111111111111010"),
    word'("111111111100110"),
    word'("111111111101110"),
    word'("111111111110100"),
    word'("111111111110111"),
    word'("111111111111010"),
    word'("111111111111100"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111101011101101"),
    word'("001111001001100"),
    word'("011010100011101"),
    word'("000001101110001"),
    word'("000100000000010"),
    word'("010101011100000"),
    word'("101011011111000"),
    word'("000000010011111"),
    word'("010001100100101"),
    word'("011110111001101"),
    word'("101000110001001"),
    word'("101111110101001"),
    word'("110100110101110"),
    word'("111000010100001"),
    word'("111010101101010"),
    word'("111100011001111"),
    word'("111101100000010"),
    word'("111110010100101"),
    word'("111110110101000"),
    word'("111111001111101"),
    word'("111111011111101"),
    word'("111111101001011"),
    word'("111111110000001"),
    word'("111111110110010"),
    word'("111111111001010"),
    word'("111111111001111"),
    word'("111111111101001"),
    word'("111111111111010"),
    word'("111111111100110"),
    word'("111111111101110"),
    word'("111111111110100"),
    word'("111111111110111"),
    word'("111111111111010"),
    word'("111111111111100"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("110000001111111"),
    word'("110111111110001"),
    word'("000011100011110"),
    word'("010011001100100"),
    word'("000000010111000"),
    word'("000110101000010"),
    word'("011001101000011"),
    word'("101111110000110"),
    word'("000100000000101"),
    word'("010100011101111"),
    word'("100001000101101"),
    word'("101010010110010"),
    word'("110000111110011"),
    word'("110101100110111"),
    word'("111000110110010"),
    word'("111011000101010"),
    word'("111100101011010"),
    word'("111101101111010"),
    word'("111110011100001"),
    word'("111110111011100"),
    word'("111111010011000"),
    word'("111111100000101"),
    word'("111111101000110"),
    word'("111111110010100"),
    word'("111111110111111"),
    word'("111111111010010"),
    word'("111111111010101"),
    word'("111111111101101"),
    word'("111111111111101"),
    word'("111111111101000"),
    word'("111111111101111"),
    word'("111111111110101"),
    word'("111111111111000"),
    word'("111111111111010"),
    word'("111111111111100"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("110000001111111"),
    word'("110111111110001"),
    word'("000011100011110"),
    word'("010011001100100"),
    word'("000000010111000"),
    word'("000110101000010"),
    word'("011001101000011"),
    word'("101111110000110"),
    word'("000100000000101"),
    word'("010100011101111"),
    word'("100001000101101"),
    word'("101010010110010"),
    word'("110000111110011"),
    word'("110101100110111"),
    word'("111000110110010"),
    word'("111011000101010"),
    word'("111100101011010"),
    word'("111101101111010"),
    word'("111110011100001"),
    word'("111110111011100"),
    word'("111111010011000"),
    word'("111111100000101"),
    word'("111111101000110"),
    word'("111111110010100"),
    word'("111111110111111"),
    word'("111111111010010"),
    word'("111111111010101"),
    word'("111111111101101"),
    word'("111111111111101"),
    word'("111111111101000"),
    word'("111111111101111"),
    word'("111111111110101"),
    word'("111111111111000"),
    word'("111111111111010"),
    word'("111111111111100"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("110110101100000"),
    word'("111100110000010"),
    word'("101011000000100"),
    word'("110010100001001"),
    word'("001010001000111"),
    word'("000000001100010"),
    word'("001011101000001"),
    word'("100000010110001"),
    word'("110110010000110"),
    word'("001001011011100"),
    word'("011000101111001"),
    word'("100100001100000"),
    word'("101100100100100"),
    word'("110010100010110"),
    word'("110110101101100"),
    word'("111001101000101"),
    word'("111011101001101"),
    word'("111101000010011"),
    word'("111101111111010"),
    word'("111110100101111"),
    word'("111111000010100"),
    word'("111111010101010"),
    word'("111111100011100"),
    word'("111111101101100"),
    word'("111111110001110"),
    word'("111111110110001"),
    word'("111111111011110"),
    word'("111111111011101"),
    word'("111111111110010"),
    word'("111111111100001"),
    word'("111111111101011"),
    word'("111111111110001"),
    word'("111111111110110"),
    word'("111111111111001"),
    word'("111111111111011"),
    word'("111111111111100"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("110110101100000"),
    word'("111100110000010"),
    word'("101011000000100"),
    word'("110010100001001"),
    word'("001010001000111"),
    word'("000000001100010"),
    word'("001011101000001"),
    word'("100000010110001"),
    word'("110110010000110"),
    word'("001001011011100"),
    word'("011000101111001"),
    word'("100100001100000"),
    word'("101100100100100"),
    word'("110010100010110"),
    word'("110110101101100"),
    word'("111001101000101"),
    word'("111011101001101"),
    word'("111101000010011"),
    word'("111101111111010"),
    word'("111110100101111"),
    word'("111111000010100"),
    word'("111111010101010"),
    word'("111111100011100"),
    word'("111111101101100"),
    word'("111111110001110"),
    word'("111111110110001"),
    word'("111111111011110"),
    word'("111111111011101"),
    word'("111111111110010"),
    word'("111111111100001"),
    word'("111111111101011"),
    word'("111111111110001"),
    word'("111111111110110"),
    word'("111111111111001"),
    word'("111111111111011"),
    word'("111111111111100"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("000101101100000"),
    word'("011010100010010"),
    word'("111111010000100"),
    word'("010101111101110"),
    word'("011111010100101"),
    word'("000010111100010"),
    word'("000010110000100"),
    word'("010011000101111"),
    word'("101000111110101"),
    word'("111110000111000"),
    word'("001111110100101"),
    word'("011101100101110"),
    word'("100111110001101"),
    word'("101111001010101"),
    word'("110100010100010"),
    word'("110111111100101"),
    word'("111010011111100"),
    word'("111100001110001"),
    word'("111101011010100"),
    word'("111110001110111"),
    word'("111110110010011"),
    word'("111111001011011"),
    word'("111111011100100"),
    word'("111111100111010"),
    word'("111111101110110"),
    word'("111111110101011"),
    word'("111111111000100"),
    word'("111111111001100"),
    word'("111111111100110"),
    word'("111111111111001"),
    word'("111111111100101"),
    word'("111111111101101"),
    word'("111111111110011"),
    word'("111111111110111"),
    word'("111111111111010"),
    word'("111111111111100"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("000101101100000"),
    word'("011010100010010"),
    word'("111111010000100"),
    word'("010101111101110"),
    word'("011111010100101"),
    word'("000010111100010"),
    word'("000010110000100"),
    word'("010011000101111"),
    word'("101000111110101"),
    word'("111110000111000"),
    word'("001111110100101"),
    word'("011101100101110"),
    word'("100111110001101"),
    word'("101111001010101"),
    word'("110100010100010"),
    word'("110111111100101"),
    word'("111010011111100"),
    word'("111100001110001"),
    word'("111101011010100"),
    word'("111110001110111"),
    word'("111110110010011"),
    word'("111111001011011"),
    word'("111111011100100"),
    word'("111111100111010"),
    word'("111111101110110"),
    word'("111111110101011"),
    word'("111111111000100"),
    word'("111111111001100"),
    word'("111111111100110"),
    word'("111111111111001"),
    word'("111111111100101"),
    word'("111111111101101"),
    word'("111111111110011"),
    word'("111111111110111"),
    word'("111111111111010"),
    word'("111111111111100"),
    word'("111111111111101"),
    word'("111111111111110"),
    word'("111111111111110"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111"),
    word'("111111111111111")
  );
BEGIN

  -- Reading ROM
  PROCESS(addr)
    VARIABLE idx_addr : INTEGER;
  BEGIN
    idx_addr := conv_integer(unsigned(addr(9 DOWNTO 0)));
    IF idx_addr >= 0 AND idx_addr < 960 THEN
      data_out <= mem(idx_addr); --spyglass disable W122 // CAT-35158
    ELSE
      data_out <= (OTHERS => '0');
    END IF;
  END PROCESS;

END v1;



--------> ./rtl_dutmgc_rom_37_960_13_1.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    2024.1_2/1117371 Production Release
--  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
-- 
--  Generated by:   dr655@ecelinux-16.ece.cornell.edu
--  Generated date: Thu Nov 28 23:23:20 2024
-- ----------------------------------------------------------------------

-- 
LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


PACKAGE dutmgc_rom_37_960_13_1_pkg IS 
  COMPONENT dutmgc_rom_37_960_13_1
    PORT (
      addr : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
    );
  END COMPONENT;
END dutmgc_rom_37_960_13_1_pkg;

PACKAGE BODY dutmgc_rom_37_960_13_1_pkg IS
END dutmgc_rom_37_960_13_1_pkg;

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


USE work.dutmgc_rom_37_960_13_1_pkg.all;
LIBRARY std;

USE std.textio.all;
USE ieee.std_logic_textio.all;

ENTITY dutmgc_rom_37_960_13_1 IS
    PORT (
      addr : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
    );
END dutmgc_rom_37_960_13_1;

ARCHITECTURE v1 OF dutmgc_rom_37_960_13_1 IS
  -- Start of SIF_NL_VHDL::nhl_rom_body
  -- Constants for ROM dimensions
  CONSTANT n_width    : INTEGER := 13;
  CONSTANT n_size     : INTEGER := 960;
  CONSTANT n_addr_w   : INTEGER := 10;
  CONSTANT n_inreg    : INTEGER := 0;
  CONSTANT n_outreg   : INTEGER := 0;
  -- Define data types for ROM storage;
  SUBTYPE  word  IS std_logic_vector((n_width)-1 DOWNTO 0);
  TYPE     lookup_table IS ARRAY (0 to n_size-1) of word;

  SIGNAL mem : lookup_table := lookup_table'(
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("0000000000000"),
    word'("1011101101010"),
    word'("1110000010100"),
    word'("0000100110011"),
    word'("0100010000110"),
    word'("1001010010111"),
    word'("1111110101110"),
    word'("0111110011000"),
    word'("0001000001110"),
    word'("1011010111011"),
    word'("0110101001010"),
    word'("0010101101101"),
    word'("1111011110000"),
    word'("1100110001101"),
    word'("1010100011001"),
    word'("1000101101100"),
    word'("0111001100100"),
    word'("0101111100000"),
    word'("0100111001101"),
    word'("0100000010111"),
    word'("0011010101110"),
    word'("0010110000011"),
    word'("0010010001100"),
    word'("0001111000001"),
    word'("0001100011001"),
    word'("0001010001111"),
    word'("0001000011100"),
    word'("0000110111110"),
    word'("0000101110000"),
    word'("0000100110000"),
    word'("0000011111011"),
    word'("0000011001111"),
    word'("0000010101010"),
    word'("0000010001101"),
    word'("0000001110100"),
    word'("0000001100000"),
    word'("0000001001111"),
    word'("0000001000001"),
    word'("0000000110110"),
    word'("0000000101100"),
    word'("0000000100100"),
    word'("0000000011110"),
    word'("0000000011001"),
    word'("0000000010100"),
    word'("0000000010001"),
    word'("0000000001110"),
    word'("0000000001011"),
    word'("0000000001001"),
    word'("0000000000111"),
    word'("1011101101010"),
    word'("1110000010100"),
    word'("0000100110011"),
    word'("0100010000110"),
    word'("1001010010111"),
    word'("1111110101110"),
    word'("0111110011000"),
    word'("0001000001110"),
    word'("1011010111011"),
    word'("0110101001010"),
    word'("0010101101101"),
    word'("1111011110000"),
    word'("1100110001101"),
    word'("1010100011001"),
    word'("1000101101100"),
    word'("0111001100100"),
    word'("0101111100000"),
    word'("0100111001101"),
    word'("0100000010111"),
    word'("0011010101110"),
    word'("0010110000011"),
    word'("0010010001100"),
    word'("0001111000001"),
    word'("0001100011001"),
    word'("0001010001111"),
    word'("0001000011100"),
    word'("0000110111110"),
    word'("0000101110000"),
    word'("0000100110000"),
    word'("0000011111011"),
    word'("0000011001111"),
    word'("0000010101010"),
    word'("0000010001101"),
    word'("0000001110100"),
    word'("0000001100000"),
    word'("0000001001111"),
    word'("0000001000001"),
    word'("0000000110110"),
    word'("0000000101100"),
    word'("0000000100100"),
    word'("0000000011110"),
    word'("0000000011001"),
    word'("0000000010100"),
    word'("0000000010001"),
    word'("0000000001110"),
    word'("0000000001011"),
    word'("0000000001001"),
    word'("0000000000111"),
    word'("0100011000111"),
    word'("1111100110000"),
    word'("1101001110100"),
    word'("0011011111011"),
    word'("0110011110001"),
    word'("1000101111110"),
    word'("1011101001101"),
    word'("1111110100011"),
    word'("0101011101110"),
    word'("1100100100111"),
    word'("0101000001101"),
    word'("1110101101101"),
    word'("1001011011000"),
    word'("0101000001110"),
    word'("0001011000100"),
    word'("1110010111100"),
    word'("1011110111011"),
    word'("1001110010111"),
    word'("1000000101101"),
    word'("0110101011100"),
    word'("0101100000111"),
    word'("0100100011001"),
    word'("0011110000011"),
    word'("0011000110011"),
    word'("0010100011110"),
    word'("0010000111001"),
    word'("0001101111100"),
    word'("0001011100000"),
    word'("0001001100000"),
    word'("0000111110110"),
    word'("0000110011110"),
    word'("0000101010101"),
    word'("0000100011010"),
    word'("0000011101001"),
    word'("0000011000000"),
    word'("0000010011110"),
    word'("0000010000011"),
    word'("0000001101100"),
    word'("0000001011001"),
    word'("0000001001001"),
    word'("0000000111100"),
    word'("0000000110010"),
    word'("0000000101001"),
    word'("0000000100010"),
    word'("0000000011100"),
    word'("0000000010111"),
    word'("0000000010011"),
    word'("0000000001111"),
    word'("0100011000111"),
    word'("1111100110000"),
    word'("1101001110100"),
    word'("0011011111011"),
    word'("0110011110001"),
    word'("1000101111110"),
    word'("1011101001101"),
    word'("1111110100011"),
    word'("0101011101110"),
    word'("1100100100111"),
    word'("0101000001101"),
    word'("1110101101101"),
    word'("1001011011000"),
    word'("0101000001110"),
    word'("0001011000100"),
    word'("1110010111100"),
    word'("1011110111011"),
    word'("1001110010111"),
    word'("1000000101101"),
    word'("0110101011100"),
    word'("0101100000111"),
    word'("0100100011001"),
    word'("0011110000011"),
    word'("0011000110011"),
    word'("0010100011110"),
    word'("0010000111001"),
    word'("0001101111100"),
    word'("0001011100000"),
    word'("0001001100000"),
    word'("0000111110110"),
    word'("0000110011110"),
    word'("0000101010101"),
    word'("0000100011010"),
    word'("0000011101001"),
    word'("0000011000000"),
    word'("0000010011110"),
    word'("0000010000011"),
    word'("0000001101100"),
    word'("0000001011001"),
    word'("0000001001001"),
    word'("0000000111100"),
    word'("0000000110010"),
    word'("0000000101001"),
    word'("0000000100010"),
    word'("0000000011100"),
    word'("0000000010111"),
    word'("0000000010011"),
    word'("0000000001111"),
    word'("0010000100000"),
    word'("1111000101011"),
    word'("0001111101110"),
    word'("1111001000010"),
    word'("1101111101111"),
    word'("0100110010100"),
    word'("1000000000010"),
    word'("1010010010011"),
    word'("1101000101111"),
    word'("0001000110100"),
    word'("0110100010101"),
    word'("1101100000010"),
    word'("0101110100010"),
    word'("1111010111010"),
    word'("1001111110010"),
    word'("0101011111101"),
    word'("0001110001000"),
    word'("1110101011001"),
    word'("1100000111110"),
    word'("1010000000111"),
    word'("1000010001001"),
    word'("0110110100101"),
    word'("0101101000101"),
    word'("0100101001101"),
    word'("0011110101110"),
    word'("0011001010110"),
    word'("0010100111011"),
    word'("0010001010001"),
    word'("0001110010000"),
    word'("0001011110001"),
    word'("0001001101101"),
    word'("0001000000000"),
    word'("0000110100111"),
    word'("0000101011101"),
    word'("0000100100000"),
    word'("0000011101110"),
    word'("0000011000100"),
    word'("0000010100010"),
    word'("0000010000101"),
    word'("0000001101110"),
    word'("0000001011011"),
    word'("0000001001011"),
    word'("0000000111110"),
    word'("0000000110011"),
    word'("0000000101010"),
    word'("0000000100010"),
    word'("0000000011100"),
    word'("0000000010111"),
    word'("0010000100000"),
    word'("1111000101011"),
    word'("0001111101110"),
    word'("1111001000010"),
    word'("1101111101111"),
    word'("0100110010100"),
    word'("1000000000010"),
    word'("1010010010011"),
    word'("1101000101111"),
    word'("0001000110100"),
    word'("0110100010101"),
    word'("1101100000010"),
    word'("0101110100010"),
    word'("1111010111010"),
    word'("1001111110010"),
    word'("0101011111101"),
    word'("0001110001000"),
    word'("1110101011001"),
    word'("1100000111110"),
    word'("1010000000111"),
    word'("1000010001001"),
    word'("0110110100101"),
    word'("0101101000101"),
    word'("0100101001101"),
    word'("0011110101110"),
    word'("0011001010110"),
    word'("0010100111011"),
    word'("0010001010001"),
    word'("0001110010000"),
    word'("0001011110001"),
    word'("0001001101101"),
    word'("0001000000000"),
    word'("0000110100111"),
    word'("0000101011101"),
    word'("0000100100000"),
    word'("0000011101110"),
    word'("0000011000100"),
    word'("0000010100010"),
    word'("0000010000101"),
    word'("0000001101110"),
    word'("0000001011011"),
    word'("0000001001011"),
    word'("0000000111110"),
    word'("0000000110011"),
    word'("0000000101010"),
    word'("0000000100010"),
    word'("0000000011100"),
    word'("0000000010111"),
    word'("1111001000010"),
    word'("1011101101011"),
    word'("0011110101110"),
    word'("0011100101111"),
    word'("1010110100000"),
    word'("1111111001111"),
    word'("1010000011000"),
    word'("1110101001000"),
    word'("0001001001111"),
    word'("0011100100101"),
    word'("0110111000101"),
    word'("1011101000011"),
    word'("0001110101011"),
    word'("1001011111001"),
    word'("0010011100011"),
    word'("1100100011011"),
    word'("0111101000010"),
    word'("0011100010000"),
    word'("0000001001001"),
    word'("1101010101111"),
    word'("1011000001001"),
    word'("1001000110000"),
    word'("0111100000101"),
    word'("0110001100110"),
    word'("0101000111101"),
    word'("0100001110011"),
    word'("0011011111001"),
    word'("0010111000001"),
    word'("0010011000000"),
    word'("0001111101100"),
    word'("0001100111100"),
    word'("0001010101011"),
    word'("0001000110100"),
    word'("0000111010010"),
    word'("0000110000000"),
    word'("0000100111101"),
    word'("0000100000110"),
    word'("0000011011000"),
    word'("0000010110010"),
    word'("0000010010011"),
    word'("0000001111001"),
    word'("0000001100100"),
    word'("0000001010010"),
    word'("0000001000100"),
    word'("0000000111000"),
    word'("0000000101110"),
    word'("0000000100110"),
    word'("0000000011111"),
    word'("1111001000010"),
    word'("1011101101011"),
    word'("0011110101110"),
    word'("0011100101111"),
    word'("1010110100000"),
    word'("1111111001111"),
    word'("1010000011000"),
    word'("1110101001000"),
    word'("0001001001111"),
    word'("0011100100101"),
    word'("0110111000101"),
    word'("1011101000011"),
    word'("0001110101011"),
    word'("1001011111001"),
    word'("0010011100011"),
    word'("1100100011011"),
    word'("0111101000010"),
    word'("0011100010000"),
    word'("0000001001001"),
    word'("1101010101111"),
    word'("1011000001001"),
    word'("1001000110000"),
    word'("0111100000101"),
    word'("0110001100110"),
    word'("0101000111101"),
    word'("0100001110011"),
    word'("0011011111001"),
    word'("0010111000001"),
    word'("0010011000000"),
    word'("0001111101100"),
    word'("0001100111100"),
    word'("0001010101011"),
    word'("0001000110100"),
    word'("0000111010010"),
    word'("0000110000000"),
    word'("0000100111101"),
    word'("0000100000110"),
    word'("0000011011000"),
    word'("0000010110010"),
    word'("0000010010011"),
    word'("0000001111001"),
    word'("0000001100100"),
    word'("0000001010010"),
    word'("0000001000100"),
    word'("0000000111000"),
    word'("0000000101110"),
    word'("0000000100110"),
    word'("0000000011111"),
    word'("0101010000011"),
    word'("0101011000101"),
    word'("1110100101000"),
    word'("1001010111100"),
    word'("1101101011010"),
    word'("1000011110101"),
    word'("1111111111100"),
    word'("1011100000001"),
    word'("0000101110011"),
    word'("0011011010000"),
    word'("0101101101001"),
    word'("1000111000100"),
    word'("1101010110100"),
    word'("0011010100111"),
    word'("1010110000011"),
    word'("0011100001100"),
    word'("1101011100001"),
    word'("1000010111001"),
    word'("0100001001100"),
    word'("0000101010010"),
    word'("1101110000110"),
    word'("1011010111001"),
    word'("1001011000101"),
    word'("0111101111111"),
    word'("0110011001100"),
    word'("0101010010000"),
    word'("0100010111000"),
    word'("0011100110010"),
    word'("0010111110001"),
    word'("0010011100111"),
    word'("0010000001100"),
    word'("0001101010110"),
    word'("0001011000010"),
    word'("0001001000110"),
    word'("0000111100000"),
    word'("0000110001100"),
    word'("0000101000111"),
    word'("0000100001110"),
    word'("0000011011111"),
    word'("0000010111000"),
    word'("0000010011000"),
    word'("0000001111101"),
    word'("0000001100111"),
    word'("0000001010101"),
    word'("0000001000110"),
    word'("0000000111010"),
    word'("0000000110000"),
    word'("0000000100111"),
    word'("0101010000011"),
    word'("0101011000101"),
    word'("1110100101000"),
    word'("1001010111100"),
    word'("1101101011010"),
    word'("1000011110101"),
    word'("1111111111100"),
    word'("1011100000001"),
    word'("0000101110011"),
    word'("0011011010000"),
    word'("0101101101001"),
    word'("1000111000100"),
    word'("1101010110100"),
    word'("0011010100111"),
    word'("1010110000011"),
    word'("0011100001100"),
    word'("1101011100001"),
    word'("1000010111001"),
    word'("0100001001100"),
    word'("0000101010010"),
    word'("1101110000110"),
    word'("1011010111001"),
    word'("1001011000101"),
    word'("0111101111111"),
    word'("0110011001100"),
    word'("0101010010000"),
    word'("0100010111000"),
    word'("0011100110010"),
    word'("0010111110001"),
    word'("0010011100111"),
    word'("0010000001100"),
    word'("0001101010110"),
    word'("0001011000010"),
    word'("0001001000110"),
    word'("0000111100000"),
    word'("0000110001100"),
    word'("0000101000111"),
    word'("0000100001110"),
    word'("0000011011111"),
    word'("0000010111000"),
    word'("0000010011000"),
    word'("0000001111101"),
    word'("0000001100111"),
    word'("0000001010101"),
    word'("0000001000110"),
    word'("0000000111010"),
    word'("0000000110000"),
    word'("0000000100111"),
    word'("1100001111000"),
    word'("0011101000011"),
    word'("1000001110110"),
    word'("0010011001001"),
    word'("1100101110001"),
    word'("1111100101110"),
    word'("1001010000000"),
    word'("1111111111111"),
    word'("1011000101010"),
    word'("0000000110101"),
    word'("0010101011110"),
    word'("0101000100001"),
    word'("1000010000100"),
    word'("1100110100010"),
    word'("0010110111100"),
    word'("1010011000010"),
    word'("0011001100000"),
    word'("1101001001111"),
    word'("1000001000101"),
    word'("0011111110000"),
    word'("0000100000000"),
    word'("1101101000000"),
    word'("1011010000100"),
    word'("1001010010111"),
    word'("0111101011010"),
    word'("0110010101100"),
    word'("0101001110110"),
    word'("0100010100010"),
    word'("0011100100001"),
    word'("0010111100010"),
    word'("0010011011011"),
    word'("0010000000001"),
    word'("0001101001111"),
    word'("0001010111011"),
    word'("0001001000001"),
    word'("0000111011100"),
    word'("0000110001001"),
    word'("0000101000100"),
    word'("0000100001011"),
    word'("0000011011101"),
    word'("0000010110110"),
    word'("0000010010110"),
    word'("0000001111100"),
    word'("0000001100110"),
    word'("0000001010100"),
    word'("0000001000101"),
    word'("0000000111001"),
    word'("0000000101111"),
    word'("1100001111000"),
    word'("0011101000011"),
    word'("1000001110110"),
    word'("0010011001001"),
    word'("1100101110001"),
    word'("1111100101110"),
    word'("1001010000000"),
    word'("1111111111111"),
    word'("1011000101010"),
    word'("0000000110101"),
    word'("0010101011110"),
    word'("0101000100001"),
    word'("1000010000100"),
    word'("1100110100010"),
    word'("0010110111100"),
    word'("1010011000010"),
    word'("0011001100000"),
    word'("1101001001111"),
    word'("1000001000101"),
    word'("0011111110000"),
    word'("0000100000000"),
    word'("1101101000000"),
    word'("1011010000100"),
    word'("1001010010111"),
    word'("0111101011010"),
    word'("0110010101100"),
    word'("0101001110110"),
    word'("0100010100010"),
    word'("0011100100001"),
    word'("0010111100010"),
    word'("0010011011011"),
    word'("0010000000001"),
    word'("0001101001111"),
    word'("0001010111011"),
    word'("0001001000001"),
    word'("0000111011100"),
    word'("0000110001001"),
    word'("0000101000100"),
    word'("0000100001011"),
    word'("0000011011101"),
    word'("0000010110110"),
    word'("0000010010110"),
    word'("0000001111100"),
    word'("0000001100110"),
    word'("0000001010100"),
    word'("0000001000101"),
    word'("0000000111001"),
    word'("0000000101111"),
    word'("0100000110000"),
    word'("0001110111100"),
    word'("0000001100101"),
    word'("0100100010110"),
    word'("0010010011100"),
    word'("1000110110010"),
    word'("0110011111010"),
    word'("1011110100110"),
    word'("1111101111111"),
    word'("1001010001000"),
    word'("1101100010101"),
    word'("0000000000000"),
    word'("0010011100010"),
    word'("0101111001001"),
    word'("1010101111101"),
    word'("0001000110100"),
    word'("1000110111001"),
    word'("0001111010000"),
    word'("1100000110001"),
    word'("0111010000110"),
    word'("0011001110110"),
    word'("1111111000101"),
    word'("1101001000010"),
    word'("1010110101111"),
    word'("1000111101000"),
    word'("0111011001000"),
    word'("0110000110100"),
    word'("0101000010010"),
    word'("0100001010001"),
    word'("0011011011101"),
    word'("0010110101010"),
    word'("0010010101100"),
    word'("0001111011100"),
    word'("0001100101111"),
    word'("0001010100001"),
    word'("0001000101011"),
    word'("0000111001010"),
    word'("0000101111010"),
    word'("0000100111000"),
    word'("0000100000001"),
    word'("0000011010100"),
    word'("0000010101111"),
    word'("0000010010001"),
    word'("0000001110111"),
    word'("0000001100010"),
    word'("0000001010001"),
    word'("0000001000011"),
    word'("0000000110111"),
    word'("0100000110000"),
    word'("0001110111100"),
    word'("0000001100101"),
    word'("0100100010110"),
    word'("0010010011100"),
    word'("1000110110010"),
    word'("0110011111010"),
    word'("1011110100110"),
    word'("1111101111111"),
    word'("1001010001000"),
    word'("1101100010101"),
    word'("0000000000000"),
    word'("0010011100010"),
    word'("0101111001001"),
    word'("1010101111101"),
    word'("0001000110100"),
    word'("1000110111001"),
    word'("0001111010000"),
    word'("1100000110001"),
    word'("0111010000110"),
    word'("0011001110110"),
    word'("1111111000101"),
    word'("1101001000010"),
    word'("1010110101111"),
    word'("1000111101000"),
    word'("0111011001000"),
    word'("0110000110100"),
    word'("0101000010010"),
    word'("0100001010001"),
    word'("0011011011101"),
    word'("0010110101010"),
    word'("0010010101100"),
    word'("0001111011100"),
    word'("0001100101111"),
    word'("0001010100001"),
    word'("0001000101011"),
    word'("0000111001010"),
    word'("0000101111010"),
    word'("0000100111000"),
    word'("0000100000001"),
    word'("0000011010100"),
    word'("0000010101111"),
    word'("0000010010001"),
    word'("0000001110111"),
    word'("0000001100010"),
    word'("0000001010001"),
    word'("0000001000011"),
    word'("0000000110111"),
    word'("1110101000110"),
    word'("1000000100010"),
    word'("0001001100111"),
    word'("0010111000000"),
    word'("1010110010011"),
    word'("1001110111010"),
    word'("1001100100010"),
    word'("1111010000111"),
    word'("1110100000100"),
    word'("1110100110100"),
    word'("0110000010111"),
    word'("1001100001111"),
    word'("1011110011011"),
    word'("1110011111101"),
    word'("0010010110010"),
    word'("0111101010111"),
    word'("1110011100100"),
    word'("0110100110111"),
    word'("0000000001111"),
    word'("1010100010100"),
    word'("0101111101000"),
    word'("0010001001000"),
    word'("1110111111110"),
    word'("1100011000110"),
    word'("1010001110110"),
    word'("1000011100100"),
    word'("0110111110010"),
    word'("0101110000011"),
    word'("0100110000001"),
    word'("0011111011000"),
    word'("0011001111001"),
    word'("0010101010111"),
    word'("0010001101001"),
    word'("0001110100100"),
    word'("0001100000001"),
    word'("0001001111010"),
    word'("0001000001100"),
    word'("0000110110000"),
    word'("0000101100101"),
    word'("0000100100110"),
    word'("0000011110011"),
    word'("0000011001000"),
    word'("0000010100101"),
    word'("0000010001000"),
    word'("0000001110000"),
    word'("0000001011101"),
    word'("0000001001100"),
    word'("0000000111111"),
    word'("1110101000110"),
    word'("1000000100010"),
    word'("0001001100111"),
    word'("0010111000000"),
    word'("1010110010011"),
    word'("1001110111010"),
    word'("1001100100010"),
    word'("1111010000111"),
    word'("1110100000100"),
    word'("1110100110100"),
    word'("0110000010111"),
    word'("1001100001111"),
    word'("1011110011011"),
    word'("1110011111101"),
    word'("0010010110010"),
    word'("0111101010111"),
    word'("1110011100100"),
    word'("0110100110111"),
    word'("0000000001111"),
    word'("1010100010100"),
    word'("0101111101000"),
    word'("0010001001000"),
    word'("1110111111110"),
    word'("1100011000110"),
    word'("1010001110110"),
    word'("1000011100100"),
    word'("0110111110010"),
    word'("0101110000011"),
    word'("0100110000001"),
    word'("0011111011000"),
    word'("0011001111001"),
    word'("0010101010111"),
    word'("0010001101001"),
    word'("0001110100100"),
    word'("0001100000001"),
    word'("0001001111010"),
    word'("0001000001100"),
    word'("0000110110000"),
    word'("0000101100101"),
    word'("0000100100110"),
    word'("0000011110011"),
    word'("0000011001000"),
    word'("0000010100101"),
    word'("0000010001000"),
    word'("0000001110000"),
    word'("0000001011101"),
    word'("0000001001100"),
    word'("0000000111111"),
    word'("0100110000000"),
    word'("0100011111101"),
    word'("1100100001000"),
    word'("0111110000111"),
    word'("0001111010010"),
    word'("1001011100110"),
    word'("0101010110101"),
    word'("1011001010110"),
    word'("0111011010101"),
    word'("1111111100010"),
    word'("1100000000110"),
    word'("0001100000101"),
    word'("0100001111111"),
    word'("0110100011111"),
    word'("1001101001010"),
    word'("1110000011111"),
    word'("0011111011100"),
    word'("1011010000001"),
    word'("0011111011101"),
    word'("1101110011001"),
    word'("1000101010100"),
    word'("0100011001000"),
    word'("0000110111000"),
    word'("1101111011011"),
    word'("1011100000011"),
    word'("1001100000000"),
    word'("0111110101111"),
    word'("0110011110011"),
    word'("0101010110001"),
    word'("0100011010011"),
    word'("0011101001000"),
    word'("0011000000010"),
    word'("0010011110111"),
    word'("0010000011001"),
    word'("0001101100001"),
    word'("0001011001010"),
    word'("0001001001110"),
    word'("0000111100110"),
    word'("0000110010001"),
    word'("0000101001011"),
    word'("0000100010001"),
    word'("0000011100001"),
    word'("0000010111010"),
    word'("0000010011001"),
    word'("0000001111111"),
    word'("0000001101000"),
    word'("0000001010110"),
    word'("0000001000111"),
    word'("0100110000000"),
    word'("0100011111101"),
    word'("1100100001000"),
    word'("0111110000111"),
    word'("0001111010010"),
    word'("1001011100110"),
    word'("0101010110101"),
    word'("1011001010110"),
    word'("0111011010101"),
    word'("1111111100010"),
    word'("1100000000110"),
    word'("0001100000101"),
    word'("0100001111111"),
    word'("0110100011111"),
    word'("1001101001010"),
    word'("1110000011111"),
    word'("0011111011100"),
    word'("1011010000001"),
    word'("0011111011101"),
    word'("1101110011001"),
    word'("1000101010100"),
    word'("0100011001000"),
    word'("0000110111000"),
    word'("1101111011011"),
    word'("1011100000011"),
    word'("1001100000000"),
    word'("0111110101111"),
    word'("0110011110011"),
    word'("0101010110001"),
    word'("0100011010011"),
    word'("0011101001000"),
    word'("0011000000010"),
    word'("0010011110111"),
    word'("0010000011001"),
    word'("0001101100001"),
    word'("0001011001010"),
    word'("0001001001110"),
    word'("0000111100110"),
    word'("0000110010001"),
    word'("0000101001011"),
    word'("0000100010001"),
    word'("0000011100001"),
    word'("0000010111010"),
    word'("0000010011001"),
    word'("0000001111111"),
    word'("0000001101000"),
    word'("0000001010110"),
    word'("0000001000111")
  );
BEGIN

  -- Reading ROM
  PROCESS(addr)
    VARIABLE idx_addr : INTEGER;
  BEGIN
    idx_addr := conv_integer(unsigned(addr(9 DOWNTO 0)));
    IF idx_addr >= 0 AND idx_addr < 960 THEN
      data_out <= mem(idx_addr); --spyglass disable W122 // CAT-35158
    ELSE
      data_out <= (OTHERS => '0');
    END IF;
  END PROCESS;

END v1;



--------> ./rtl_dutmgc_rom_38_64_8_1.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    2024.1_2/1117371 Production Release
--  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
-- 
--  Generated by:   dr655@ecelinux-16.ece.cornell.edu
--  Generated date: Thu Nov 28 23:23:20 2024
-- ----------------------------------------------------------------------

-- 
LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


PACKAGE dutmgc_rom_38_64_8_1_pkg IS 
  COMPONENT dutmgc_rom_38_64_8_1
    PORT (
      addr : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
  END COMPONENT;
END dutmgc_rom_38_64_8_1_pkg;

PACKAGE BODY dutmgc_rom_38_64_8_1_pkg IS
END dutmgc_rom_38_64_8_1_pkg;

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


USE work.dutmgc_rom_38_64_8_1_pkg.all;
LIBRARY std;

USE std.textio.all;
USE ieee.std_logic_textio.all;

ENTITY dutmgc_rom_38_64_8_1 IS
    PORT (
      addr : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END dutmgc_rom_38_64_8_1;

ARCHITECTURE v1 OF dutmgc_rom_38_64_8_1 IS
  -- Start of SIF_NL_VHDL::nhl_rom_body
  -- Constants for ROM dimensions
  CONSTANT n_width    : INTEGER := 8;
  CONSTANT n_size     : INTEGER := 64;
  CONSTANT n_addr_w   : INTEGER := 6;
  CONSTANT n_inreg    : INTEGER := 0;
  CONSTANT n_outreg   : INTEGER := 0;
  -- Define data types for ROM storage;
  SUBTYPE  word  IS std_logic_vector((n_width)-1 DOWNTO 0);
  TYPE     lookup_table IS ARRAY (0 to n_size-1) of word;

  SIGNAL mem : lookup_table := lookup_table'(
    word'("00001010"),
    word'("00100010"),
    word'("01100101"),
    word'("00010010"),
    word'("00000001"),
    word'("10101001"),
    word'("00100001"),
    word'("01011010"),
    word'("01010001"),
    word'("01000101"),
    word'("00000101"),
    word'("10010101"),
    word'("10011010"),
    word'("10001000"),
    word'("01011001"),
    word'("10001001"),
    word'("10011010"),
    word'("10101000"),
    word'("10101010"),
    word'("01100100"),
    word'("01001010"),
    word'("00000101"),
    word'("01010110"),
    word'("01010001"),
    word'("10100110"),
    word'("00101001"),
    word'("01000001"),
    word'("10011001"),
    word'("00010101"),
    word'("10101001"),
    word'("01010110"),
    word'("10100101"),
    word'("10101001"),
    word'("10000010"),
    word'("00100101"),
    word'("01010010"),
    word'("10000010"),
    word'("01010110"),
    word'("10010010"),
    word'("01001000"),
    word'("10010100"),
    word'("10010001"),
    word'("01100101"),
    word'("01010000"),
    word'("01011010"),
    word'("01100001"),
    word'("01101010"),
    word'("10100000"),
    word'("10010000"),
    word'("01010100"),
    word'("01010000"),
    word'("01010101"),
    word'("01011000"),
    word'("01001001"),
    word'("01011001"),
    word'("00000110"),
    word'("10000100"),
    word'("10100110"),
    word'("10010101"),
    word'("10000110"),
    word'("00010110"),
    word'("10101000"),
    word'("10100010"),
    word'("01001010")
  );
BEGIN

  -- Reading ROM
  PROCESS(addr)
    VARIABLE idx_addr : INTEGER;
  BEGIN
    idx_addr := conv_integer(unsigned(addr(5 DOWNTO 0)));
    data_out <= mem(idx_addr); --spyglass disable W122 // CAT-35158
  END PROCESS;

END v1;



--------> ./rtl_dutmgc_rom_39_64_8_1.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    2024.1_2/1117371 Production Release
--  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
-- 
--  Generated by:   dr655@ecelinux-16.ece.cornell.edu
--  Generated date: Thu Nov 28 23:23:20 2024
-- ----------------------------------------------------------------------

-- 
LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


PACKAGE dutmgc_rom_39_64_8_1_pkg IS 
  COMPONENT dutmgc_rom_39_64_8_1
    PORT (
      addr : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
  END COMPONENT;
END dutmgc_rom_39_64_8_1_pkg;

PACKAGE BODY dutmgc_rom_39_64_8_1_pkg IS
END dutmgc_rom_39_64_8_1_pkg;

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


USE work.dutmgc_rom_39_64_8_1_pkg.all;
LIBRARY std;

USE std.textio.all;
USE ieee.std_logic_textio.all;

ENTITY dutmgc_rom_39_64_8_1 IS
    PORT (
      addr : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END dutmgc_rom_39_64_8_1;

ARCHITECTURE v1 OF dutmgc_rom_39_64_8_1 IS
  -- Start of SIF_NL_VHDL::nhl_rom_body
  -- Constants for ROM dimensions
  CONSTANT n_width    : INTEGER := 8;
  CONSTANT n_size     : INTEGER := 64;
  CONSTANT n_addr_w   : INTEGER := 6;
  CONSTANT n_inreg    : INTEGER := 0;
  CONSTANT n_outreg   : INTEGER := 0;
  -- Define data types for ROM storage;
  SUBTYPE  word  IS std_logic_vector((n_width)-1 DOWNTO 0);
  TYPE     lookup_table IS ARRAY (0 to n_size-1) of word;

  SIGNAL mem : lookup_table := lookup_table'(
    word'("10000010"),
    word'("00011001"),
    word'("01000101"),
    word'("10101000"),
    word'("00011001"),
    word'("00001010"),
    word'("10010101"),
    word'("00010100"),
    word'("00010101"),
    word'("10010000"),
    word'("00001001"),
    word'("01100010"),
    word'("10001010"),
    word'("10010010"),
    word'("01010001"),
    word'("01101010"),
    word'("10100001"),
    word'("01100110"),
    word'("00101000"),
    word'("01010000"),
    word'("01101000"),
    word'("00100000"),
    word'("10100101"),
    word'("10100100"),
    word'("10010010"),
    word'("00000010"),
    word'("01101000"),
    word'("10010001"),
    word'("00101000"),
    word'("00011010"),
    word'("10000010"),
    word'("01011010"),
    word'("00000010"),
    word'("00001001"),
    word'("00000101"),
    word'("01000101"),
    word'("10001000"),
    word'("01100010"),
    word'("00001001"),
    word'("10010010"),
    word'("00000001"),
    word'("01101001"),
    word'("01101001"),
    word'("00100101"),
    word'("00010100"),
    word'("00001000"),
    word'("00101010"),
    word'("10011010"),
    word'("00010100"),
    word'("01101001"),
    word'("00100110"),
    word'("10010000"),
    word'("10001000"),
    word'("10010000"),
    word'("00000100"),
    word'("00010000"),
    word'("10101000"),
    word'("00011000"),
    word'("00000100"),
    word'("10010000"),
    word'("01100110"),
    word'("00011000"),
    word'("00010000"),
    word'("00010100")
  );
BEGIN

  -- Reading ROM
  PROCESS(addr)
    VARIABLE idx_addr : INTEGER;
  BEGIN
    idx_addr := conv_integer(unsigned(addr(5 DOWNTO 0)));
    data_out <= mem(idx_addr); --spyglass disable W122 // CAT-35158
  END PROCESS;

END v1;



--------> ./rtl_dutmgc_rom_40_32_19_1.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    2024.1_2/1117371 Production Release
--  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
-- 
--  Generated by:   dr655@ecelinux-16.ece.cornell.edu
--  Generated date: Thu Nov 28 23:23:20 2024
-- ----------------------------------------------------------------------

-- 
LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


PACKAGE dutmgc_rom_40_32_19_1_pkg IS 
  COMPONENT dutmgc_rom_40_32_19_1
    PORT (
      addr : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
    );
  END COMPONENT;
END dutmgc_rom_40_32_19_1_pkg;

PACKAGE BODY dutmgc_rom_40_32_19_1_pkg IS
END dutmgc_rom_40_32_19_1_pkg;

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


USE work.dutmgc_rom_40_32_19_1_pkg.all;
LIBRARY std;

USE std.textio.all;
USE ieee.std_logic_textio.all;

ENTITY dutmgc_rom_40_32_19_1 IS
    PORT (
      addr : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
    );
END dutmgc_rom_40_32_19_1;

ARCHITECTURE v1 OF dutmgc_rom_40_32_19_1 IS
  -- Start of SIF_NL_VHDL::nhl_rom_body
  -- Constants for ROM dimensions
  CONSTANT n_width    : INTEGER := 19;
  CONSTANT n_size     : INTEGER := 32;
  CONSTANT n_addr_w   : INTEGER := 5;
  CONSTANT n_inreg    : INTEGER := 0;
  CONSTANT n_outreg   : INTEGER := 0;
  -- Define data types for ROM storage;
  SUBTYPE  word  IS std_logic_vector((n_width)-1 DOWNTO 0);
  TYPE     lookup_table IS ARRAY (0 to n_size-1) of word;

  SIGNAL mem : lookup_table := lookup_table'(
    word'("0000000000101000010"),
    word'("0000001010001111110"),
    word'("1111101100100110111"),
    word'("0000001000110101000"),
    word'("1111111111101011110"),
    word'("0000001000001100101"),
    word'("1111010101010001101"),
    word'("1111110000100011001"),
    word'("0000010000001111001"),
    word'("0000000010101011100"),
    word'("0000000001111001000"),
    word'("1111101110010101111"),
    word'("1010110101101110011"),
    word'("1111000101010001000"),
    word'("0011111100000101010"),
    word'("0010100100101111011"),
    word'("0000010110011000101"),
    word'("1111111010101000111"),
    word'("0000001001001001001"),
    word'("1111111010011110110"),
    word'("1100000010011111010"),
    word'("0010000100001011101"),
    word'("0010111101010111111"),
    word'("0100000100000111010"),
    word'("0000000001100100111"),
    word'("1111111101111100110"),
    word'("0000000011011101111"),
    word'("1111100111111000010"),
    word'("1110010000011101100"),
    word'("1110011010101110011"),
    word'("0011110000011010100"),
    word'("0001000001000001000")
  );
BEGIN

  -- Reading ROM
  PROCESS(addr)
    VARIABLE idx_addr : INTEGER;
  BEGIN
    idx_addr := conv_integer(unsigned(addr(4 DOWNTO 0)));
    data_out <= mem(idx_addr); --spyglass disable W122 // CAT-35158
  END PROCESS;

END v1;



--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    2024.1_2/1117371 Production Release
--  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
-- 
--  Generated by:   dr655@ecelinux-16.ece.cornell.edu
--  Generated date: Thu Nov 28 23:23:20 2024
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_16_6_40_48_1_48_40_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_16_6_40_48_1_48_40_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
    re : OUT STD_LOGIC;
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    re_d : IN STD_LOGIC;
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_16_6_40_48_1_48_40_1_gen;

ARCHITECTURE v1 OF dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_16_6_40_48_1_48_40_1_gen
    IS
  CONSTANT PowerPro_35032 : STD_LOGIC := '1';
BEGIN
  clken <= (clken_d);
  q_d <= q;
  re <= (readA_r_ram_ir_internal_RMASK_B_d);
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_15_6_40_48_1_48_40_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_15_6_40_48_1_48_40_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
    re : OUT STD_LOGIC;
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    re_d : IN STD_LOGIC;
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_15_6_40_48_1_48_40_1_gen;

ARCHITECTURE v1 OF dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_15_6_40_48_1_48_40_1_gen
    IS
  CONSTANT PowerPro_35032 : STD_LOGIC := '1';
BEGIN
  clken <= (clken_d);
  q_d <= q;
  re <= (readA_r_ram_ir_internal_RMASK_B_d);
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_14_6_40_48_1_48_40_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_14_6_40_48_1_48_40_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
    re : OUT STD_LOGIC;
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    re_d : IN STD_LOGIC;
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_14_6_40_48_1_48_40_1_gen;

ARCHITECTURE v1 OF dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_14_6_40_48_1_48_40_1_gen
    IS
  CONSTANT PowerPro_35032 : STD_LOGIC := '1';
BEGIN
  clken <= (clken_d);
  q_d <= q;
  re <= (readA_r_ram_ir_internal_RMASK_B_d);
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    dut_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY dut_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    for_for_C_2_tr0 : IN STD_LOGIC;
    compute_sqrt_for_C_15_tr0 : IN STD_LOGIC;
    RMS_NORM_LOOP_2_C_4_tr0 : IN STD_LOGIC;
    QUANTIZE_ACTIVATION_LOOP_3_C_2_tr0 : IN STD_LOGIC;
    LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0 : IN STD_LOGIC;
    LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0 : IN STD_LOGIC;
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_63_tr0 : IN STD_LOGIC;
    RESHAPE_2D_TO_3D_LOOP_3_C_0_tr0 : IN STD_LOGIC;
    RESHAPE_2D_TO_3D_LOOP_2_C_0_tr0 : IN STD_LOGIC;
    RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0 : IN STD_LOGIC;
    RESHAPE_2D_TO_3D_LOOP_2_2_C_0_tr0 : IN STD_LOGIC;
    APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0 : IN STD_LOGIC;
    APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0 : IN STD_LOGIC;
    CACHE_UPDATE_LOOP_3_C_1_tr0 : IN STD_LOGIC;
    CACHE_UPDATE_LOOP_2_C_0_tr0 : IN STD_LOGIC;
    CACHE_UPDATE_LOOP_1_C_0_tr0 : IN STD_LOGIC;
    TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0 : IN STD_LOGIC;
    TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0 : IN STD_LOGIC;
    TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0 : IN STD_LOGIC;
    GEMM_3D_FLOAT_LOOP_4_C_3_tr0 : IN STD_LOGIC;
    GEMM_3D_FLOAT_LOOP_3_C_1_tr0 : IN STD_LOGIC;
    GEMM_3D_FLOAT_LOOP_1_C_0_tr0 : IN STD_LOGIC;
    SF_LOOP_3_C_0_tr0 : IN STD_LOGIC;
    SF_LOOP_1_C_0_tr0 : IN STD_LOGIC;
    CM_LOOP_1_C_0_tr0 : IN STD_LOGIC;
    SOFTMAX_LOOP_3_C_0_tr0 : IN STD_LOGIC;
    SOFTMAX_LOOP_4_C_2_tr0 : IN STD_LOGIC;
    SOFTMAX_LOOP_5_C_19_tr0 : IN STD_LOGIC;
    SOFTMAX_LOOP_1_C_1_tr0 : IN STD_LOGIC;
    GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0 : IN STD_LOGIC;
    GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0 : IN STD_LOGIC;
    GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0 : IN STD_LOGIC;
    ATTN_2D_LOOP_3_C_0_tr0 : IN STD_LOGIC;
    ATTN_2D_LOOP_2_C_0_tr0 : IN STD_LOGIC;
    RMS_NORM_LOOP_1_2_C_2_tr0 : IN STD_LOGIC;
    compute_sqrt_1_for_C_15_tr0 : IN STD_LOGIC;
    RMS_NORM_LOOP_2_2_C_4_tr0 : IN STD_LOGIC;
    QUANTIZE_ACTIVATION_LOOP_3_1_C_2_tr0 : IN STD_LOGIC;
    LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0 : IN STD_LOGIC;
    LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0 : IN STD_LOGIC;
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31_tr0 : IN STD_LOGIC;
    for_1_for_C_1_tr0 : IN STD_LOGIC
  );
END dut_core_core_fsm;

ARCHITECTURE v1 OF dut_core_core_fsm IS
  -- FSM State Type Declaration for dut_core_core_fsm_1
  TYPE dut_core_core_fsm_1_ST IS (main_C_0, for_for_C_0, for_for_C_1, for_for_C_2,
      main_C_1, compute_sqrt_for_C_0, compute_sqrt_for_C_1, compute_sqrt_for_C_2,
      compute_sqrt_for_C_3, compute_sqrt_for_C_4, compute_sqrt_for_C_5, compute_sqrt_for_C_6,
      compute_sqrt_for_C_7, compute_sqrt_for_C_8, compute_sqrt_for_C_9, compute_sqrt_for_C_10,
      compute_sqrt_for_C_11, compute_sqrt_for_C_12, compute_sqrt_for_C_13, compute_sqrt_for_C_14,
      compute_sqrt_for_C_15, main_C_2, main_C_3, main_C_4, main_C_5, main_C_6, main_C_7,
      main_C_8, main_C_9, main_C_10, main_C_11, main_C_12, main_C_13, main_C_14,
      main_C_15, main_C_16, main_C_17, main_C_18, main_C_19, main_C_20, main_C_21,
      main_C_22, main_C_23, main_C_24, main_C_25, main_C_26, main_C_27, main_C_28,
      main_C_29, main_C_30, main_C_31, main_C_32, main_C_33, RMS_NORM_LOOP_2_C_0,
      RMS_NORM_LOOP_2_C_1, RMS_NORM_LOOP_2_C_2, RMS_NORM_LOOP_2_C_3, RMS_NORM_LOOP_2_C_4,
      main_C_34, main_C_35, main_C_36, main_C_37, main_C_38, main_C_39, main_C_40,
      main_C_41, main_C_42, main_C_43, main_C_44, main_C_45, main_C_46, main_C_47,
      main_C_48, QUANTIZE_ACTIVATION_LOOP_3_C_0, QUANTIZE_ACTIVATION_LOOP_3_C_1,
      QUANTIZE_ACTIVATION_LOOP_3_C_2, LINEAR_FORWARD_NO_MUL_LOOP_3_C_0, LINEAR_FORWARD_NO_MUL_LOOP_4_C_0,
      LINEAR_FORWARD_NO_MUL_LOOP_3_C_1, LINEAR_FORWARD_NO_MUL_LOOP_2_C_0, LINEAR_FORWARD_NO_MUL_LOOP_2_C_1,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_2, LINEAR_FORWARD_NO_MUL_LOOP_2_C_3, LINEAR_FORWARD_NO_MUL_LOOP_2_C_4,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_5, LINEAR_FORWARD_NO_MUL_LOOP_2_C_6, LINEAR_FORWARD_NO_MUL_LOOP_2_C_7,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_8, LINEAR_FORWARD_NO_MUL_LOOP_2_C_9, LINEAR_FORWARD_NO_MUL_LOOP_2_C_10,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_11, LINEAR_FORWARD_NO_MUL_LOOP_2_C_12, LINEAR_FORWARD_NO_MUL_LOOP_2_C_13,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_14, LINEAR_FORWARD_NO_MUL_LOOP_2_C_15, LINEAR_FORWARD_NO_MUL_LOOP_2_C_16,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_17, LINEAR_FORWARD_NO_MUL_LOOP_2_C_18, LINEAR_FORWARD_NO_MUL_LOOP_2_C_19,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_20, LINEAR_FORWARD_NO_MUL_LOOP_2_C_21, LINEAR_FORWARD_NO_MUL_LOOP_2_C_22,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_23, LINEAR_FORWARD_NO_MUL_LOOP_2_C_24, LINEAR_FORWARD_NO_MUL_LOOP_2_C_25,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_26, LINEAR_FORWARD_NO_MUL_LOOP_2_C_27, LINEAR_FORWARD_NO_MUL_LOOP_2_C_28,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_29, LINEAR_FORWARD_NO_MUL_LOOP_2_C_30, LINEAR_FORWARD_NO_MUL_LOOP_2_C_31,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_32, LINEAR_FORWARD_NO_MUL_LOOP_2_C_33, LINEAR_FORWARD_NO_MUL_LOOP_2_C_34,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_35, LINEAR_FORWARD_NO_MUL_LOOP_2_C_36, LINEAR_FORWARD_NO_MUL_LOOP_2_C_37,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_38, LINEAR_FORWARD_NO_MUL_LOOP_2_C_39, LINEAR_FORWARD_NO_MUL_LOOP_2_C_40,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_41, LINEAR_FORWARD_NO_MUL_LOOP_2_C_42, LINEAR_FORWARD_NO_MUL_LOOP_2_C_43,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_44, LINEAR_FORWARD_NO_MUL_LOOP_2_C_45, LINEAR_FORWARD_NO_MUL_LOOP_2_C_46,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_47, LINEAR_FORWARD_NO_MUL_LOOP_2_C_48, LINEAR_FORWARD_NO_MUL_LOOP_2_C_49,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_50, LINEAR_FORWARD_NO_MUL_LOOP_2_C_51, LINEAR_FORWARD_NO_MUL_LOOP_2_C_52,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_53, LINEAR_FORWARD_NO_MUL_LOOP_2_C_54, LINEAR_FORWARD_NO_MUL_LOOP_2_C_55,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_56, LINEAR_FORWARD_NO_MUL_LOOP_2_C_57, LINEAR_FORWARD_NO_MUL_LOOP_2_C_58,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_59, LINEAR_FORWARD_NO_MUL_LOOP_2_C_60, LINEAR_FORWARD_NO_MUL_LOOP_2_C_61,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_62, LINEAR_FORWARD_NO_MUL_LOOP_2_C_63, RESHAPE_2D_TO_3D_LOOP_3_C_0,
      RESHAPE_2D_TO_3D_LOOP_2_C_0, RESHAPE_2D_TO_3D_LOOP_3_2_C_0, RESHAPE_2D_TO_3D_LOOP_2_2_C_0,
      APPLY_ROTARY_POS_EMB_LOOP_6_C_0, APPLY_ROTARY_POS_EMB_LOOP_6_C_1, APPLY_ROTARY_POS_EMB_LOOP_6_C_2,
      APPLY_ROTARY_POS_EMB_LOOP_4_C_0, CACHE_UPDATE_LOOP_3_C_0, CACHE_UPDATE_LOOP_3_C_1,
      CACHE_UPDATE_LOOP_2_C_0, CACHE_UPDATE_LOOP_1_C_0, TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_0,
      TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_1, TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2, TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0,
      TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0, GEMM_3D_FLOAT_LOOP_3_C_0, GEMM_3D_FLOAT_LOOP_4_C_0,
      GEMM_3D_FLOAT_LOOP_4_C_1, GEMM_3D_FLOAT_LOOP_4_C_2, GEMM_3D_FLOAT_LOOP_4_C_3,
      GEMM_3D_FLOAT_LOOP_3_C_1, GEMM_3D_FLOAT_LOOP_1_C_0, SF_LOOP_3_C_0, SF_LOOP_1_C_0,
      CM_LOOP_1_C_0, SOFTMAX_LOOP_1_C_0, SOFTMAX_LOOP_3_C_0, SOFTMAX_LOOP_4_C_0,
      SOFTMAX_LOOP_4_C_1, SOFTMAX_LOOP_4_C_2, SOFTMAX_LOOP_5_C_0, SOFTMAX_LOOP_5_C_1,
      SOFTMAX_LOOP_5_C_2, SOFTMAX_LOOP_5_C_3, SOFTMAX_LOOP_5_C_4, SOFTMAX_LOOP_5_C_5,
      SOFTMAX_LOOP_5_C_6, SOFTMAX_LOOP_5_C_7, SOFTMAX_LOOP_5_C_8, SOFTMAX_LOOP_5_C_9,
      SOFTMAX_LOOP_5_C_10, SOFTMAX_LOOP_5_C_11, SOFTMAX_LOOP_5_C_12, SOFTMAX_LOOP_5_C_13,
      SOFTMAX_LOOP_5_C_14, SOFTMAX_LOOP_5_C_15, SOFTMAX_LOOP_5_C_16, SOFTMAX_LOOP_5_C_17,
      SOFTMAX_LOOP_5_C_18, SOFTMAX_LOOP_5_C_19, SOFTMAX_LOOP_1_C_1, GEMM_3D_FLOAT_LOOP_3_1_C_0,
      GEMM_3D_FLOAT_LOOP_4_1_C_0, GEMM_3D_FLOAT_LOOP_4_1_C_1, GEMM_3D_FLOAT_LOOP_4_1_C_2,
      GEMM_3D_FLOAT_LOOP_4_1_C_3, GEMM_3D_FLOAT_LOOP_3_1_C_1, GEMM_3D_FLOAT_LOOP_1_1_C_0,
      ATTN_2D_LOOP_3_C_0, ATTN_2D_LOOP_2_C_0, RMS_NORM_LOOP_1_2_C_0, RMS_NORM_LOOP_1_2_C_1,
      RMS_NORM_LOOP_1_2_C_2, main_C_49, compute_sqrt_1_for_C_0, compute_sqrt_1_for_C_1,
      compute_sqrt_1_for_C_2, compute_sqrt_1_for_C_3, compute_sqrt_1_for_C_4, compute_sqrt_1_for_C_5,
      compute_sqrt_1_for_C_6, compute_sqrt_1_for_C_7, compute_sqrt_1_for_C_8, compute_sqrt_1_for_C_9,
      compute_sqrt_1_for_C_10, compute_sqrt_1_for_C_11, compute_sqrt_1_for_C_12,
      compute_sqrt_1_for_C_13, compute_sqrt_1_for_C_14, compute_sqrt_1_for_C_15,
      main_C_50, main_C_51, main_C_52, main_C_53, main_C_54, main_C_55, main_C_56,
      main_C_57, main_C_58, main_C_59, main_C_60, main_C_61, main_C_62, main_C_63,
      main_C_64, main_C_65, main_C_66, main_C_67, main_C_68, RMS_NORM_LOOP_2_2_C_0,
      RMS_NORM_LOOP_2_2_C_1, RMS_NORM_LOOP_2_2_C_2, RMS_NORM_LOOP_2_2_C_3, RMS_NORM_LOOP_2_2_C_4,
      main_C_69, main_C_70, main_C_71, main_C_72, main_C_73, main_C_74, main_C_75,
      main_C_76, main_C_77, main_C_78, main_C_79, main_C_80, main_C_81, main_C_82,
      main_C_83, main_C_84, main_C_85, main_C_86, main_C_87, main_C_88, main_C_89,
      main_C_90, main_C_91, main_C_92, main_C_93, main_C_94, main_C_95, main_C_96,
      main_C_97, main_C_98, main_C_99, main_C_100, QUANTIZE_ACTIVATION_LOOP_3_1_C_0,
      QUANTIZE_ACTIVATION_LOOP_3_1_C_1, QUANTIZE_ACTIVATION_LOOP_3_1_C_2, LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_0,
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0, LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_0,
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_1, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_2, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_3,
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_4, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_5, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_6,
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_7, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_8, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_9,
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_10, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_11, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_12,
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_13, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_14, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_15,
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_16, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_17, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_18,
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_19, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_20, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_21,
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_22, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_23, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_24,
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_25, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_26, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_27,
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_28, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_29, LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_30,
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31, for_1_for_C_0, for_1_for_C_1);

  SIGNAL state_var : dut_core_core_fsm_1_ST;
  SIGNAL state_var_NS : dut_core_core_fsm_1_ST;

BEGIN
  dut_core_core_fsm_1 : PROCESS (for_for_C_2_tr0, compute_sqrt_for_C_15_tr0, RMS_NORM_LOOP_2_C_4_tr0,
      QUANTIZE_ACTIVATION_LOOP_3_C_2_tr0, LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0, LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_63_tr0, RESHAPE_2D_TO_3D_LOOP_3_C_0_tr0, RESHAPE_2D_TO_3D_LOOP_2_C_0_tr0,
      RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0, RESHAPE_2D_TO_3D_LOOP_2_2_C_0_tr0, APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0,
      APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0, CACHE_UPDATE_LOOP_3_C_1_tr0, CACHE_UPDATE_LOOP_2_C_0_tr0,
      CACHE_UPDATE_LOOP_1_C_0_tr0, TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0, TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0,
      TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0, GEMM_3D_FLOAT_LOOP_4_C_3_tr0, GEMM_3D_FLOAT_LOOP_3_C_1_tr0,
      GEMM_3D_FLOAT_LOOP_1_C_0_tr0, SF_LOOP_3_C_0_tr0, SF_LOOP_1_C_0_tr0, CM_LOOP_1_C_0_tr0,
      SOFTMAX_LOOP_3_C_0_tr0, SOFTMAX_LOOP_4_C_2_tr0, SOFTMAX_LOOP_5_C_19_tr0, SOFTMAX_LOOP_1_C_1_tr0,
      GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0, GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0, GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0,
      ATTN_2D_LOOP_3_C_0_tr0, ATTN_2D_LOOP_2_C_0_tr0, RMS_NORM_LOOP_1_2_C_2_tr0,
      compute_sqrt_1_for_C_15_tr0, RMS_NORM_LOOP_2_2_C_4_tr0, QUANTIZE_ACTIVATION_LOOP_3_1_C_2_tr0,
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0, LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0,
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31_tr0, for_1_for_C_1_tr0, state_var)
  BEGIN
    CASE state_var IS
      WHEN for_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000001");
        state_var_NS <= for_for_C_1;
      WHEN for_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000010");
        state_var_NS <= for_for_C_2;
      WHEN for_for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000011");
        IF ( for_for_C_2_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSE
          state_var_NS <= for_for_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000100");
        state_var_NS <= compute_sqrt_for_C_0;
      WHEN compute_sqrt_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000101");
        state_var_NS <= compute_sqrt_for_C_1;
      WHEN compute_sqrt_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000110");
        state_var_NS <= compute_sqrt_for_C_2;
      WHEN compute_sqrt_for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000111");
        state_var_NS <= compute_sqrt_for_C_3;
      WHEN compute_sqrt_for_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001000");
        state_var_NS <= compute_sqrt_for_C_4;
      WHEN compute_sqrt_for_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001001");
        state_var_NS <= compute_sqrt_for_C_5;
      WHEN compute_sqrt_for_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001010");
        state_var_NS <= compute_sqrt_for_C_6;
      WHEN compute_sqrt_for_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001011");
        state_var_NS <= compute_sqrt_for_C_7;
      WHEN compute_sqrt_for_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001100");
        state_var_NS <= compute_sqrt_for_C_8;
      WHEN compute_sqrt_for_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001101");
        state_var_NS <= compute_sqrt_for_C_9;
      WHEN compute_sqrt_for_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001110");
        state_var_NS <= compute_sqrt_for_C_10;
      WHEN compute_sqrt_for_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001111");
        state_var_NS <= compute_sqrt_for_C_11;
      WHEN compute_sqrt_for_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010000");
        state_var_NS <= compute_sqrt_for_C_12;
      WHEN compute_sqrt_for_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010001");
        state_var_NS <= compute_sqrt_for_C_13;
      WHEN compute_sqrt_for_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010010");
        state_var_NS <= compute_sqrt_for_C_14;
      WHEN compute_sqrt_for_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010011");
        state_var_NS <= compute_sqrt_for_C_15;
      WHEN compute_sqrt_for_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010100");
        IF ( compute_sqrt_for_C_15_tr0 = '1' ) THEN
          state_var_NS <= main_C_2;
        ELSE
          state_var_NS <= compute_sqrt_for_C_0;
        END IF;
      WHEN main_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010101");
        state_var_NS <= main_C_3;
      WHEN main_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010110");
        state_var_NS <= main_C_4;
      WHEN main_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010111");
        state_var_NS <= main_C_5;
      WHEN main_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011000");
        state_var_NS <= main_C_6;
      WHEN main_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011001");
        state_var_NS <= main_C_7;
      WHEN main_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011010");
        state_var_NS <= main_C_8;
      WHEN main_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011011");
        state_var_NS <= main_C_9;
      WHEN main_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011100");
        state_var_NS <= main_C_10;
      WHEN main_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011101");
        state_var_NS <= main_C_11;
      WHEN main_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011110");
        state_var_NS <= main_C_12;
      WHEN main_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011111");
        state_var_NS <= main_C_13;
      WHEN main_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100000");
        state_var_NS <= main_C_14;
      WHEN main_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100001");
        state_var_NS <= main_C_15;
      WHEN main_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100010");
        state_var_NS <= main_C_16;
      WHEN main_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100011");
        state_var_NS <= main_C_17;
      WHEN main_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100100");
        state_var_NS <= main_C_18;
      WHEN main_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100101");
        state_var_NS <= main_C_19;
      WHEN main_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100110");
        state_var_NS <= main_C_20;
      WHEN main_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100111");
        state_var_NS <= main_C_21;
      WHEN main_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101000");
        state_var_NS <= main_C_22;
      WHEN main_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101001");
        state_var_NS <= main_C_23;
      WHEN main_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101010");
        state_var_NS <= main_C_24;
      WHEN main_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101011");
        state_var_NS <= main_C_25;
      WHEN main_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101100");
        state_var_NS <= main_C_26;
      WHEN main_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101101");
        state_var_NS <= main_C_27;
      WHEN main_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101110");
        state_var_NS <= main_C_28;
      WHEN main_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101111");
        state_var_NS <= main_C_29;
      WHEN main_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110000");
        state_var_NS <= main_C_30;
      WHEN main_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110001");
        state_var_NS <= main_C_31;
      WHEN main_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110010");
        state_var_NS <= main_C_32;
      WHEN main_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110011");
        state_var_NS <= main_C_33;
      WHEN main_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110100");
        state_var_NS <= RMS_NORM_LOOP_2_C_0;
      WHEN RMS_NORM_LOOP_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110101");
        state_var_NS <= RMS_NORM_LOOP_2_C_1;
      WHEN RMS_NORM_LOOP_2_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110110");
        state_var_NS <= RMS_NORM_LOOP_2_C_2;
      WHEN RMS_NORM_LOOP_2_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110111");
        state_var_NS <= RMS_NORM_LOOP_2_C_3;
      WHEN RMS_NORM_LOOP_2_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111000");
        state_var_NS <= RMS_NORM_LOOP_2_C_4;
      WHEN RMS_NORM_LOOP_2_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111001");
        IF ( RMS_NORM_LOOP_2_C_4_tr0 = '1' ) THEN
          state_var_NS <= main_C_34;
        ELSE
          state_var_NS <= RMS_NORM_LOOP_2_C_0;
        END IF;
      WHEN main_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111010");
        state_var_NS <= main_C_35;
      WHEN main_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111011");
        state_var_NS <= main_C_36;
      WHEN main_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111100");
        state_var_NS <= main_C_37;
      WHEN main_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111101");
        state_var_NS <= main_C_38;
      WHEN main_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111110");
        state_var_NS <= main_C_39;
      WHEN main_C_39 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111111");
        state_var_NS <= main_C_40;
      WHEN main_C_40 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000000");
        state_var_NS <= main_C_41;
      WHEN main_C_41 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000001");
        state_var_NS <= main_C_42;
      WHEN main_C_42 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000010");
        state_var_NS <= main_C_43;
      WHEN main_C_43 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000011");
        state_var_NS <= main_C_44;
      WHEN main_C_44 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000100");
        state_var_NS <= main_C_45;
      WHEN main_C_45 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000101");
        state_var_NS <= main_C_46;
      WHEN main_C_46 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000110");
        state_var_NS <= main_C_47;
      WHEN main_C_47 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000111");
        state_var_NS <= main_C_48;
      WHEN main_C_48 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001000");
        state_var_NS <= QUANTIZE_ACTIVATION_LOOP_3_C_0;
      WHEN QUANTIZE_ACTIVATION_LOOP_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001001");
        state_var_NS <= QUANTIZE_ACTIVATION_LOOP_3_C_1;
      WHEN QUANTIZE_ACTIVATION_LOOP_3_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001010");
        state_var_NS <= QUANTIZE_ACTIVATION_LOOP_3_C_2;
      WHEN QUANTIZE_ACTIVATION_LOOP_3_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001011");
        IF ( QUANTIZE_ACTIVATION_LOOP_3_C_2_tr0 = '1' ) THEN
          state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_3_C_0;
        ELSE
          state_var_NS <= QUANTIZE_ACTIVATION_LOOP_3_C_0;
        END IF;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001100");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_4_C_0;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_4_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001101");
        IF ( LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0 = '1' ) THEN
          state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_3_C_1;
        ELSE
          state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_4_C_0;
        END IF;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_3_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001110");
        IF ( LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0 = '1' ) THEN
          state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_0;
        ELSE
          state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_3_C_0;
        END IF;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001111");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_1;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010000");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_2;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010001");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_3;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010010");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_4;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010011");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_5;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010100");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_6;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010101");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_7;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010110");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_8;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010111");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_9;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011000");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_10;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011001");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_11;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011010");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_12;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011011");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_13;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011100");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_14;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011101");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_15;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011110");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_16;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011111");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_17;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100000");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_18;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100001");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_19;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100010");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_20;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100011");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_21;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100100");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_22;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100101");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_23;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100110");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_24;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100111");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_25;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101000");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_26;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101001");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_27;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101010");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_28;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101011");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_29;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101100");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_30;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101101");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_31;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101110");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_32;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101111");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_33;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110000");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_34;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110001");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_35;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110010");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_36;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110011");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_37;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110100");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_38;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110101");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_39;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_39 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110110");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_40;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_40 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110111");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_41;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_41 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111000");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_42;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_42 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111001");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_43;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_43 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111010");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_44;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_44 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111011");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_45;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_45 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111100");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_46;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_46 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111101");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_47;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_47 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111110");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_48;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_48 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111111");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_49;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_49 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000000");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_50;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_50 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000001");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_51;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_51 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000010");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_52;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_52 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000011");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_53;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_53 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000100");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_54;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_54 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000101");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_55;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_55 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000110");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_56;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_56 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000111");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_57;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_57 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001000");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_58;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_58 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001001");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_59;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_59 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001010");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_60;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_60 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001011");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_61;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_61 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001100");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_62;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_62 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001101");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_C_63;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_C_63 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001110");
        IF ( LINEAR_FORWARD_NO_MUL_LOOP_2_C_63_tr0 = '1' ) THEN
          state_var_NS <= RESHAPE_2D_TO_3D_LOOP_3_C_0;
        ELSE
          state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_3_C_0;
        END IF;
      WHEN RESHAPE_2D_TO_3D_LOOP_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001111");
        IF ( RESHAPE_2D_TO_3D_LOOP_3_C_0_tr0 = '1' ) THEN
          state_var_NS <= RESHAPE_2D_TO_3D_LOOP_2_C_0;
        ELSE
          state_var_NS <= RESHAPE_2D_TO_3D_LOOP_3_C_0;
        END IF;
      WHEN RESHAPE_2D_TO_3D_LOOP_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010000");
        IF ( RESHAPE_2D_TO_3D_LOOP_2_C_0_tr0 = '1' ) THEN
          state_var_NS <= RESHAPE_2D_TO_3D_LOOP_3_2_C_0;
        ELSE
          state_var_NS <= RESHAPE_2D_TO_3D_LOOP_3_C_0;
        END IF;
      WHEN RESHAPE_2D_TO_3D_LOOP_3_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010001");
        IF ( RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0 = '1' ) THEN
          state_var_NS <= RESHAPE_2D_TO_3D_LOOP_2_2_C_0;
        ELSE
          state_var_NS <= RESHAPE_2D_TO_3D_LOOP_3_2_C_0;
        END IF;
      WHEN RESHAPE_2D_TO_3D_LOOP_2_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010010");
        IF ( RESHAPE_2D_TO_3D_LOOP_2_2_C_0_tr0 = '1' ) THEN
          state_var_NS <= APPLY_ROTARY_POS_EMB_LOOP_6_C_0;
        ELSE
          state_var_NS <= RESHAPE_2D_TO_3D_LOOP_3_2_C_0;
        END IF;
      WHEN APPLY_ROTARY_POS_EMB_LOOP_6_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010011");
        state_var_NS <= APPLY_ROTARY_POS_EMB_LOOP_6_C_1;
      WHEN APPLY_ROTARY_POS_EMB_LOOP_6_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010100");
        state_var_NS <= APPLY_ROTARY_POS_EMB_LOOP_6_C_2;
      WHEN APPLY_ROTARY_POS_EMB_LOOP_6_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010101");
        IF ( APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0 = '1' ) THEN
          state_var_NS <= APPLY_ROTARY_POS_EMB_LOOP_4_C_0;
        ELSE
          state_var_NS <= APPLY_ROTARY_POS_EMB_LOOP_6_C_0;
        END IF;
      WHEN APPLY_ROTARY_POS_EMB_LOOP_4_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010110");
        IF ( APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0 = '1' ) THEN
          state_var_NS <= CACHE_UPDATE_LOOP_3_C_0;
        ELSE
          state_var_NS <= APPLY_ROTARY_POS_EMB_LOOP_6_C_0;
        END IF;
      WHEN CACHE_UPDATE_LOOP_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010111");
        state_var_NS <= CACHE_UPDATE_LOOP_3_C_1;
      WHEN CACHE_UPDATE_LOOP_3_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011000");
        IF ( CACHE_UPDATE_LOOP_3_C_1_tr0 = '1' ) THEN
          state_var_NS <= CACHE_UPDATE_LOOP_2_C_0;
        ELSE
          state_var_NS <= CACHE_UPDATE_LOOP_3_C_0;
        END IF;
      WHEN CACHE_UPDATE_LOOP_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011001");
        IF ( CACHE_UPDATE_LOOP_2_C_0_tr0 = '1' ) THEN
          state_var_NS <= CACHE_UPDATE_LOOP_1_C_0;
        ELSE
          state_var_NS <= CACHE_UPDATE_LOOP_3_C_0;
        END IF;
      WHEN CACHE_UPDATE_LOOP_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011010");
        IF ( CACHE_UPDATE_LOOP_1_C_0_tr0 = '1' ) THEN
          state_var_NS <= TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_0;
        ELSE
          state_var_NS <= CACHE_UPDATE_LOOP_3_C_0;
        END IF;
      WHEN TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011011");
        state_var_NS <= TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_1;
      WHEN TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011100");
        state_var_NS <= TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2;
      WHEN TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011101");
        IF ( TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0 = '1' ) THEN
          state_var_NS <= TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0;
        ELSE
          state_var_NS <= TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_0;
        END IF;
      WHEN TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011110");
        IF ( TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0 = '1' ) THEN
          state_var_NS <= TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0;
        ELSE
          state_var_NS <= TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_0;
        END IF;
      WHEN TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011111");
        IF ( TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0 = '1' ) THEN
          state_var_NS <= GEMM_3D_FLOAT_LOOP_3_C_0;
        ELSE
          state_var_NS <= TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_0;
        END IF;
      WHEN GEMM_3D_FLOAT_LOOP_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100000");
        state_var_NS <= GEMM_3D_FLOAT_LOOP_4_C_0;
      WHEN GEMM_3D_FLOAT_LOOP_4_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100001");
        state_var_NS <= GEMM_3D_FLOAT_LOOP_4_C_1;
      WHEN GEMM_3D_FLOAT_LOOP_4_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100010");
        state_var_NS <= GEMM_3D_FLOAT_LOOP_4_C_2;
      WHEN GEMM_3D_FLOAT_LOOP_4_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100011");
        state_var_NS <= GEMM_3D_FLOAT_LOOP_4_C_3;
      WHEN GEMM_3D_FLOAT_LOOP_4_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100100");
        IF ( GEMM_3D_FLOAT_LOOP_4_C_3_tr0 = '1' ) THEN
          state_var_NS <= GEMM_3D_FLOAT_LOOP_3_C_1;
        ELSE
          state_var_NS <= GEMM_3D_FLOAT_LOOP_4_C_0;
        END IF;
      WHEN GEMM_3D_FLOAT_LOOP_3_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100101");
        IF ( GEMM_3D_FLOAT_LOOP_3_C_1_tr0 = '1' ) THEN
          state_var_NS <= GEMM_3D_FLOAT_LOOP_1_C_0;
        ELSE
          state_var_NS <= GEMM_3D_FLOAT_LOOP_3_C_0;
        END IF;
      WHEN GEMM_3D_FLOAT_LOOP_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100110");
        IF ( GEMM_3D_FLOAT_LOOP_1_C_0_tr0 = '1' ) THEN
          state_var_NS <= SF_LOOP_3_C_0;
        ELSE
          state_var_NS <= GEMM_3D_FLOAT_LOOP_3_C_0;
        END IF;
      WHEN SF_LOOP_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100111");
        IF ( SF_LOOP_3_C_0_tr0 = '1' ) THEN
          state_var_NS <= SF_LOOP_1_C_0;
        ELSE
          state_var_NS <= SF_LOOP_3_C_0;
        END IF;
      WHEN SF_LOOP_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101000");
        IF ( SF_LOOP_1_C_0_tr0 = '1' ) THEN
          state_var_NS <= CM_LOOP_1_C_0;
        ELSE
          state_var_NS <= SF_LOOP_3_C_0;
        END IF;
      WHEN CM_LOOP_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101001");
        IF ( CM_LOOP_1_C_0_tr0 = '1' ) THEN
          state_var_NS <= SOFTMAX_LOOP_1_C_0;
        ELSE
          state_var_NS <= CM_LOOP_1_C_0;
        END IF;
      WHEN SOFTMAX_LOOP_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101010");
        state_var_NS <= SOFTMAX_LOOP_3_C_0;
      WHEN SOFTMAX_LOOP_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101011");
        IF ( SOFTMAX_LOOP_3_C_0_tr0 = '1' ) THEN
          state_var_NS <= SOFTMAX_LOOP_4_C_0;
        ELSE
          state_var_NS <= SOFTMAX_LOOP_3_C_0;
        END IF;
      WHEN SOFTMAX_LOOP_4_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101100");
        state_var_NS <= SOFTMAX_LOOP_4_C_1;
      WHEN SOFTMAX_LOOP_4_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101101");
        state_var_NS <= SOFTMAX_LOOP_4_C_2;
      WHEN SOFTMAX_LOOP_4_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101110");
        IF ( SOFTMAX_LOOP_4_C_2_tr0 = '1' ) THEN
          state_var_NS <= SOFTMAX_LOOP_5_C_0;
        ELSE
          state_var_NS <= SOFTMAX_LOOP_4_C_0;
        END IF;
      WHEN SOFTMAX_LOOP_5_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101111");
        state_var_NS <= SOFTMAX_LOOP_5_C_1;
      WHEN SOFTMAX_LOOP_5_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110000");
        state_var_NS <= SOFTMAX_LOOP_5_C_2;
      WHEN SOFTMAX_LOOP_5_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110001");
        state_var_NS <= SOFTMAX_LOOP_5_C_3;
      WHEN SOFTMAX_LOOP_5_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110010");
        state_var_NS <= SOFTMAX_LOOP_5_C_4;
      WHEN SOFTMAX_LOOP_5_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110011");
        state_var_NS <= SOFTMAX_LOOP_5_C_5;
      WHEN SOFTMAX_LOOP_5_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110100");
        state_var_NS <= SOFTMAX_LOOP_5_C_6;
      WHEN SOFTMAX_LOOP_5_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110101");
        state_var_NS <= SOFTMAX_LOOP_5_C_7;
      WHEN SOFTMAX_LOOP_5_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110110");
        state_var_NS <= SOFTMAX_LOOP_5_C_8;
      WHEN SOFTMAX_LOOP_5_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110111");
        state_var_NS <= SOFTMAX_LOOP_5_C_9;
      WHEN SOFTMAX_LOOP_5_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111000");
        state_var_NS <= SOFTMAX_LOOP_5_C_10;
      WHEN SOFTMAX_LOOP_5_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111001");
        state_var_NS <= SOFTMAX_LOOP_5_C_11;
      WHEN SOFTMAX_LOOP_5_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111010");
        state_var_NS <= SOFTMAX_LOOP_5_C_12;
      WHEN SOFTMAX_LOOP_5_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111011");
        state_var_NS <= SOFTMAX_LOOP_5_C_13;
      WHEN SOFTMAX_LOOP_5_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111100");
        state_var_NS <= SOFTMAX_LOOP_5_C_14;
      WHEN SOFTMAX_LOOP_5_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111101");
        state_var_NS <= SOFTMAX_LOOP_5_C_15;
      WHEN SOFTMAX_LOOP_5_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111110");
        state_var_NS <= SOFTMAX_LOOP_5_C_16;
      WHEN SOFTMAX_LOOP_5_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111111");
        state_var_NS <= SOFTMAX_LOOP_5_C_17;
      WHEN SOFTMAX_LOOP_5_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000000");
        state_var_NS <= SOFTMAX_LOOP_5_C_18;
      WHEN SOFTMAX_LOOP_5_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000001");
        state_var_NS <= SOFTMAX_LOOP_5_C_19;
      WHEN SOFTMAX_LOOP_5_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000010");
        IF ( SOFTMAX_LOOP_5_C_19_tr0 = '1' ) THEN
          state_var_NS <= SOFTMAX_LOOP_1_C_1;
        ELSE
          state_var_NS <= SOFTMAX_LOOP_5_C_0;
        END IF;
      WHEN SOFTMAX_LOOP_1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000011");
        IF ( SOFTMAX_LOOP_1_C_1_tr0 = '1' ) THEN
          state_var_NS <= GEMM_3D_FLOAT_LOOP_3_1_C_0;
        ELSE
          state_var_NS <= SOFTMAX_LOOP_1_C_0;
        END IF;
      WHEN GEMM_3D_FLOAT_LOOP_3_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000100");
        state_var_NS <= GEMM_3D_FLOAT_LOOP_4_1_C_0;
      WHEN GEMM_3D_FLOAT_LOOP_4_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000101");
        state_var_NS <= GEMM_3D_FLOAT_LOOP_4_1_C_1;
      WHEN GEMM_3D_FLOAT_LOOP_4_1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000110");
        state_var_NS <= GEMM_3D_FLOAT_LOOP_4_1_C_2;
      WHEN GEMM_3D_FLOAT_LOOP_4_1_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000111");
        state_var_NS <= GEMM_3D_FLOAT_LOOP_4_1_C_3;
      WHEN GEMM_3D_FLOAT_LOOP_4_1_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001000");
        IF ( GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0 = '1' ) THEN
          state_var_NS <= GEMM_3D_FLOAT_LOOP_3_1_C_1;
        ELSE
          state_var_NS <= GEMM_3D_FLOAT_LOOP_4_1_C_0;
        END IF;
      WHEN GEMM_3D_FLOAT_LOOP_3_1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001001");
        IF ( GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0 = '1' ) THEN
          state_var_NS <= GEMM_3D_FLOAT_LOOP_1_1_C_0;
        ELSE
          state_var_NS <= GEMM_3D_FLOAT_LOOP_3_1_C_0;
        END IF;
      WHEN GEMM_3D_FLOAT_LOOP_1_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001010");
        IF ( GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0 = '1' ) THEN
          state_var_NS <= ATTN_2D_LOOP_3_C_0;
        ELSE
          state_var_NS <= GEMM_3D_FLOAT_LOOP_3_1_C_0;
        END IF;
      WHEN ATTN_2D_LOOP_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001011");
        IF ( ATTN_2D_LOOP_3_C_0_tr0 = '1' ) THEN
          state_var_NS <= ATTN_2D_LOOP_2_C_0;
        ELSE
          state_var_NS <= ATTN_2D_LOOP_3_C_0;
        END IF;
      WHEN ATTN_2D_LOOP_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001100");
        IF ( ATTN_2D_LOOP_2_C_0_tr0 = '1' ) THEN
          state_var_NS <= RMS_NORM_LOOP_1_2_C_0;
        ELSE
          state_var_NS <= ATTN_2D_LOOP_3_C_0;
        END IF;
      WHEN RMS_NORM_LOOP_1_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001101");
        state_var_NS <= RMS_NORM_LOOP_1_2_C_1;
      WHEN RMS_NORM_LOOP_1_2_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001110");
        state_var_NS <= RMS_NORM_LOOP_1_2_C_2;
      WHEN RMS_NORM_LOOP_1_2_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001111");
        IF ( RMS_NORM_LOOP_1_2_C_2_tr0 = '1' ) THEN
          state_var_NS <= main_C_49;
        ELSE
          state_var_NS <= RMS_NORM_LOOP_1_2_C_0;
        END IF;
      WHEN main_C_49 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010000");
        state_var_NS <= compute_sqrt_1_for_C_0;
      WHEN compute_sqrt_1_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010001");
        state_var_NS <= compute_sqrt_1_for_C_1;
      WHEN compute_sqrt_1_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010010");
        state_var_NS <= compute_sqrt_1_for_C_2;
      WHEN compute_sqrt_1_for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010011");
        state_var_NS <= compute_sqrt_1_for_C_3;
      WHEN compute_sqrt_1_for_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010100");
        state_var_NS <= compute_sqrt_1_for_C_4;
      WHEN compute_sqrt_1_for_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010101");
        state_var_NS <= compute_sqrt_1_for_C_5;
      WHEN compute_sqrt_1_for_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010110");
        state_var_NS <= compute_sqrt_1_for_C_6;
      WHEN compute_sqrt_1_for_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010111");
        state_var_NS <= compute_sqrt_1_for_C_7;
      WHEN compute_sqrt_1_for_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011000");
        state_var_NS <= compute_sqrt_1_for_C_8;
      WHEN compute_sqrt_1_for_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011001");
        state_var_NS <= compute_sqrt_1_for_C_9;
      WHEN compute_sqrt_1_for_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011010");
        state_var_NS <= compute_sqrt_1_for_C_10;
      WHEN compute_sqrt_1_for_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011011");
        state_var_NS <= compute_sqrt_1_for_C_11;
      WHEN compute_sqrt_1_for_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011100");
        state_var_NS <= compute_sqrt_1_for_C_12;
      WHEN compute_sqrt_1_for_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011101");
        state_var_NS <= compute_sqrt_1_for_C_13;
      WHEN compute_sqrt_1_for_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011110");
        state_var_NS <= compute_sqrt_1_for_C_14;
      WHEN compute_sqrt_1_for_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011111");
        state_var_NS <= compute_sqrt_1_for_C_15;
      WHEN compute_sqrt_1_for_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100000");
        IF ( compute_sqrt_1_for_C_15_tr0 = '1' ) THEN
          state_var_NS <= main_C_50;
        ELSE
          state_var_NS <= compute_sqrt_1_for_C_0;
        END IF;
      WHEN main_C_50 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100001");
        state_var_NS <= main_C_51;
      WHEN main_C_51 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100010");
        state_var_NS <= main_C_52;
      WHEN main_C_52 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100011");
        state_var_NS <= main_C_53;
      WHEN main_C_53 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100100");
        state_var_NS <= main_C_54;
      WHEN main_C_54 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100101");
        state_var_NS <= main_C_55;
      WHEN main_C_55 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100110");
        state_var_NS <= main_C_56;
      WHEN main_C_56 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100111");
        state_var_NS <= main_C_57;
      WHEN main_C_57 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101000");
        state_var_NS <= main_C_58;
      WHEN main_C_58 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101001");
        state_var_NS <= main_C_59;
      WHEN main_C_59 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101010");
        state_var_NS <= main_C_60;
      WHEN main_C_60 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101011");
        state_var_NS <= main_C_61;
      WHEN main_C_61 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101100");
        state_var_NS <= main_C_62;
      WHEN main_C_62 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101101");
        state_var_NS <= main_C_63;
      WHEN main_C_63 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101110");
        state_var_NS <= main_C_64;
      WHEN main_C_64 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101111");
        state_var_NS <= main_C_65;
      WHEN main_C_65 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110000");
        state_var_NS <= main_C_66;
      WHEN main_C_66 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110001");
        state_var_NS <= main_C_67;
      WHEN main_C_67 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110010");
        state_var_NS <= main_C_68;
      WHEN main_C_68 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110011");
        state_var_NS <= RMS_NORM_LOOP_2_2_C_0;
      WHEN RMS_NORM_LOOP_2_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110100");
        state_var_NS <= RMS_NORM_LOOP_2_2_C_1;
      WHEN RMS_NORM_LOOP_2_2_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110101");
        state_var_NS <= RMS_NORM_LOOP_2_2_C_2;
      WHEN RMS_NORM_LOOP_2_2_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110110");
        state_var_NS <= RMS_NORM_LOOP_2_2_C_3;
      WHEN RMS_NORM_LOOP_2_2_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110111");
        state_var_NS <= RMS_NORM_LOOP_2_2_C_4;
      WHEN RMS_NORM_LOOP_2_2_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111000");
        IF ( RMS_NORM_LOOP_2_2_C_4_tr0 = '1' ) THEN
          state_var_NS <= main_C_69;
        ELSE
          state_var_NS <= RMS_NORM_LOOP_2_2_C_0;
        END IF;
      WHEN main_C_69 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111001");
        state_var_NS <= main_C_70;
      WHEN main_C_70 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111010");
        state_var_NS <= main_C_71;
      WHEN main_C_71 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111011");
        state_var_NS <= main_C_72;
      WHEN main_C_72 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111100");
        state_var_NS <= main_C_73;
      WHEN main_C_73 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111101");
        state_var_NS <= main_C_74;
      WHEN main_C_74 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111110");
        state_var_NS <= main_C_75;
      WHEN main_C_75 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111111");
        state_var_NS <= main_C_76;
      WHEN main_C_76 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000000");
        state_var_NS <= main_C_77;
      WHEN main_C_77 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000001");
        state_var_NS <= main_C_78;
      WHEN main_C_78 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000010");
        state_var_NS <= main_C_79;
      WHEN main_C_79 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000011");
        state_var_NS <= main_C_80;
      WHEN main_C_80 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000100");
        state_var_NS <= main_C_81;
      WHEN main_C_81 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000101");
        state_var_NS <= main_C_82;
      WHEN main_C_82 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000110");
        state_var_NS <= main_C_83;
      WHEN main_C_83 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000111");
        state_var_NS <= main_C_84;
      WHEN main_C_84 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001000");
        state_var_NS <= main_C_85;
      WHEN main_C_85 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001001");
        state_var_NS <= main_C_86;
      WHEN main_C_86 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001010");
        state_var_NS <= main_C_87;
      WHEN main_C_87 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001011");
        state_var_NS <= main_C_88;
      WHEN main_C_88 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001100");
        state_var_NS <= main_C_89;
      WHEN main_C_89 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001101");
        state_var_NS <= main_C_90;
      WHEN main_C_90 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001110");
        state_var_NS <= main_C_91;
      WHEN main_C_91 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001111");
        state_var_NS <= main_C_92;
      WHEN main_C_92 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010000");
        state_var_NS <= main_C_93;
      WHEN main_C_93 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010001");
        state_var_NS <= main_C_94;
      WHEN main_C_94 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010010");
        state_var_NS <= main_C_95;
      WHEN main_C_95 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010011");
        state_var_NS <= main_C_96;
      WHEN main_C_96 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010100");
        state_var_NS <= main_C_97;
      WHEN main_C_97 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010101");
        state_var_NS <= main_C_98;
      WHEN main_C_98 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010110");
        state_var_NS <= main_C_99;
      WHEN main_C_99 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010111");
        state_var_NS <= main_C_100;
      WHEN main_C_100 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011000");
        state_var_NS <= QUANTIZE_ACTIVATION_LOOP_3_1_C_0;
      WHEN QUANTIZE_ACTIVATION_LOOP_3_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011001");
        state_var_NS <= QUANTIZE_ACTIVATION_LOOP_3_1_C_1;
      WHEN QUANTIZE_ACTIVATION_LOOP_3_1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011010");
        state_var_NS <= QUANTIZE_ACTIVATION_LOOP_3_1_C_2;
      WHEN QUANTIZE_ACTIVATION_LOOP_3_1_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011011");
        IF ( QUANTIZE_ACTIVATION_LOOP_3_1_C_2_tr0 = '1' ) THEN
          state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_0;
        ELSE
          state_var_NS <= QUANTIZE_ACTIVATION_LOOP_3_1_C_0;
        END IF;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011100");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011101");
        IF ( LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0 = '1' ) THEN
          state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1;
        ELSE
          state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0;
        END IF;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011110");
        IF ( LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0 = '1' ) THEN
          state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_0;
        ELSE
          state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_0;
        END IF;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011111");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_1;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100000");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_2;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100001");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_3;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100010");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_4;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100011");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_5;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100100");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_6;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100101");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_7;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100110");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_8;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100111");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_9;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101000");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_10;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101001");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_11;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101010");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_12;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101011");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_13;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101100");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_14;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101101");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_15;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101110");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_16;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101111");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_17;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110000");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_18;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110001");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_19;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110010");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_20;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110011");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_21;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110100");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_22;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110101");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_23;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110110");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_24;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110111");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_25;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111000");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_26;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111001");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_27;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111010");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_28;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111011");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_29;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111100");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_30;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111101");
        state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31;
      WHEN LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111110");
        IF ( LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31_tr0 = '1' ) THEN
          state_var_NS <= for_1_for_C_0;
        ELSE
          state_var_NS <= LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_0;
        END IF;
      WHEN for_1_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111111");
        state_var_NS <= for_1_for_C_1;
      WHEN for_1_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101000000");
        IF ( for_1_for_C_1_tr0 = '1' ) THEN
          state_var_NS <= main_C_0;
        ELSE
          state_var_NS <= for_1_for_C_0;
        END IF;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000000");
        state_var_NS <= for_for_C_0;
    END CASE;
  END PROCESS dut_core_core_fsm_1;

  dut_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        IF ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 = '1' ) THEN
          state_var <= state_var_NS;
        END IF;
      END IF;
    END IF;
  END PROCESS dut_core_core_fsm_1_REG;

END v1;

-- ------------------------------------------------------------------
--  Design Unit:    dut_core_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY dut_core_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    rms_norm_16_div_cmp_z : IN STD_LOGIC_VECTOR (71 DOWNTO 0);
    core_wen1 : IN STD_LOGIC;
    rms_norm_16_div_cmp_z_oreg : OUT STD_LOGIC_VECTOR (39 DOWNTO 0)
  );
END dut_core_wait_dp;

ARCHITECTURE v1 OF dut_core_wait_dp IS
  -- Interconnect Declarations
  SIGNAL rms_norm_16_div_cmp_z_oreg_pconst_39_0 : STD_LOGIC_VECTOR (39 DOWNTO 0);

BEGIN
  rms_norm_16_div_cmp_z_oreg <= rms_norm_16_div_cmp_z_oreg_pconst_39_0;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        rms_norm_16_div_cmp_z_oreg_pconst_39_0 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( core_wen1 = '1' ) THEN
        rms_norm_16_div_cmp_z_oreg_pconst_39_0 <= rms_norm_16_div_cmp_z(39 DOWNTO
            0);
      END IF;
    END IF;
  END PROCESS;
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    dut_core_staller
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY dut_core_staller IS
  PORT(
    en : IN STD_LOGIC;
    core_wen1 : OUT STD_LOGIC;
    strm_in_rsci_wen_comp : IN STD_LOGIC;
    strm_out_rsci_wen_comp : IN STD_LOGIC;
    attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 : OUT STD_LOGIC
  );
END dut_core_staller;

ARCHITECTURE v1 OF dut_core_staller IS
  -- Output Reader Declarations
  SIGNAL core_wen1_drv : STD_LOGIC;

BEGIN
  -- Output Reader Assignments
  core_wen1 <= core_wen1_drv;

  attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 <= core_wen1_drv AND en;
  core_wen1_drv <= strm_in_rsci_wen_comp AND strm_out_rsci_wen_comp;
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    dut_core_strm_out_rsci_strm_out_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY dut_core_strm_out_rsci_strm_out_wait_ctrl IS
  PORT(
    strm_out_rsci_iswt0 : IN STD_LOGIC;
    strm_out_rsci_biwt : OUT STD_LOGIC;
    strm_out_rsci_irdy : IN STD_LOGIC
  );
END dut_core_strm_out_rsci_strm_out_wait_ctrl;

ARCHITECTURE v1 OF dut_core_strm_out_rsci_strm_out_wait_ctrl IS
  CONSTANT PowerPro_35032 : STD_LOGIC := '1';
BEGIN
  strm_out_rsci_biwt <= strm_out_rsci_iswt0 AND strm_out_rsci_irdy;
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    dut_core_strm_in_rsci_strm_in_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY dut_core_strm_in_rsci_strm_in_wait_ctrl IS
  PORT(
    strm_in_rsci_iswt0 : IN STD_LOGIC;
    strm_in_rsci_biwt : OUT STD_LOGIC;
    strm_in_rsci_ivld : IN STD_LOGIC
  );
END dut_core_strm_in_rsci_strm_in_wait_ctrl;

ARCHITECTURE v1 OF dut_core_strm_in_rsci_strm_in_wait_ctrl IS
  CONSTANT PowerPro_35032 : STD_LOGIC := '1';
BEGIN
  strm_in_rsci_biwt <= strm_in_rsci_iswt0 AND strm_in_rsci_ivld;
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    dut_core_strm_out_rsci
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY dut_core_strm_out_rsci IS
  PORT(
    strm_out_rsc_dat : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    strm_out_rsc_vld : OUT STD_LOGIC;
    strm_out_rsc_rdy : IN STD_LOGIC;
    strm_out_rsci_oswt : IN STD_LOGIC;
    strm_out_rsci_wen_comp : OUT STD_LOGIC;
    strm_out_rsci_idat : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END dut_core_strm_out_rsci;

ARCHITECTURE v1 OF dut_core_strm_out_rsci IS
  -- Interconnect Declarations
  SIGNAL strm_out_rsci_biwt : STD_LOGIC;
  SIGNAL strm_out_rsci_irdy : STD_LOGIC;

  SIGNAL strm_out_rsci_idat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL strm_out_rsci_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT dut_core_strm_out_rsci_strm_out_wait_ctrl
    PORT(
      strm_out_rsci_iswt0 : IN STD_LOGIC;
      strm_out_rsci_biwt : OUT STD_LOGIC;
      strm_out_rsci_irdy : IN STD_LOGIC
    );
  END COMPONENT;
BEGIN
  strm_out_rsci : work.ccs_out_wait_pkg_v1.ccs_out_wait_v1
    GENERIC MAP(
      rscid => 2,
      width => 32
      )
    PORT MAP(
      irdy => strm_out_rsci_irdy,
      ivld => strm_out_rsci_oswt,
      idat => strm_out_rsci_idat_1,
      rdy => strm_out_rsc_rdy,
      vld => strm_out_rsc_vld,
      dat => strm_out_rsci_dat
    );
  strm_out_rsci_idat_1 <= (strm_out_rsci_idat(31 DOWNTO 2)) & STD_LOGIC_VECTOR'(
      "00");
  strm_out_rsc_dat <= strm_out_rsci_dat;

  dut_core_strm_out_rsci_strm_out_wait_ctrl_inst : dut_core_strm_out_rsci_strm_out_wait_ctrl
    PORT MAP(
      strm_out_rsci_iswt0 => strm_out_rsci_oswt,
      strm_out_rsci_biwt => strm_out_rsci_biwt,
      strm_out_rsci_irdy => strm_out_rsci_irdy
    );
  strm_out_rsci_wen_comp <= (NOT strm_out_rsci_oswt) OR strm_out_rsci_biwt;
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    dut_core_strm_in_rsci
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY dut_core_strm_in_rsci IS
  PORT(
    strm_in_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    strm_in_rsc_vld : IN STD_LOGIC;
    strm_in_rsc_rdy : OUT STD_LOGIC;
    strm_in_rsci_oswt : IN STD_LOGIC;
    strm_in_rsci_wen_comp : OUT STD_LOGIC;
    strm_in_rsci_idat_mxwt : OUT STD_LOGIC_VECTOR (29 DOWNTO 0)
  );
END dut_core_strm_in_rsci;

ARCHITECTURE v1 OF dut_core_strm_in_rsci IS
  -- Interconnect Declarations
  SIGNAL strm_in_rsci_biwt : STD_LOGIC;
  SIGNAL strm_in_rsci_ivld : STD_LOGIC;
  SIGNAL strm_in_rsci_idat : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL strm_in_rsci_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL strm_in_rsci_idat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT dut_core_strm_in_rsci_strm_in_wait_ctrl
    PORT(
      strm_in_rsci_iswt0 : IN STD_LOGIC;
      strm_in_rsci_biwt : OUT STD_LOGIC;
      strm_in_rsci_ivld : IN STD_LOGIC
    );
  END COMPONENT;
BEGIN
  strm_in_rsci : work.ccs_in_wait_pkg_v1.ccs_in_wait_v1
    GENERIC MAP(
      rscid => 1,
      width => 32
      )
    PORT MAP(
      rdy => strm_in_rsc_rdy,
      vld => strm_in_rsc_vld,
      dat => strm_in_rsci_dat,
      irdy => strm_in_rsci_oswt,
      ivld => strm_in_rsci_ivld,
      idat => strm_in_rsci_idat_1
    );
  strm_in_rsci_dat <= strm_in_rsc_dat;
  strm_in_rsci_idat <= strm_in_rsci_idat_1;

  dut_core_strm_in_rsci_strm_in_wait_ctrl_inst : dut_core_strm_in_rsci_strm_in_wait_ctrl
    PORT MAP(
      strm_in_rsci_iswt0 => strm_in_rsci_oswt,
      strm_in_rsci_biwt => strm_in_rsci_biwt,
      strm_in_rsci_ivld => strm_in_rsci_ivld
    );
  strm_in_rsci_idat_mxwt <= strm_in_rsci_idat(31 DOWNTO 2);
  strm_in_rsci_wen_comp <= (NOT strm_in_rsci_oswt) OR strm_in_rsci_biwt;
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    dut_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY dut_core IS
  PORT(
    clk : IN STD_LOGIC;
    en : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    strm_in_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    strm_in_rsc_vld : IN STD_LOGIC;
    strm_in_rsc_rdy : OUT STD_LOGIC;
    strm_out_rsc_dat : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    strm_out_rsc_vld : OUT STD_LOGIC;
    strm_out_rsc_rdy : IN STD_LOGIC;
    attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d : OUT STD_LOGIC;
    attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d : OUT STD_LOGIC_VECTOR (39 DOWNTO
        0);
    attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d : OUT STD_LOGIC_VECTOR (5 DOWNTO
        0);
    attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d : OUT STD_LOGIC_VECTOR (5 DOWNTO
        0);
    attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d : OUT STD_LOGIC_VECTOR (39 DOWNTO
        0);
    attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d : IN STD_LOGIC_VECTOR (39 DOWNTO
        0);
    attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d : OUT STD_LOGIC_VECTOR (5 DOWNTO
        0);
    attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d : OUT STD_LOGIC_VECTOR (5 DOWNTO
        0);
    attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d : IN STD_LOGIC_VECTOR (39
        DOWNTO 0);
    attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d : OUT STD_LOGIC_VECTOR
        (5 DOWNTO 0);
    attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d : OUT STD_LOGIC_VECTOR
        (5 DOWNTO 0);
    rms_norm_16_div_cmp_a : OUT STD_LOGIC_VECTOR (71 DOWNTO 0);
    rms_norm_16_div_cmp_b : OUT STD_LOGIC_VECTOR (60 DOWNTO 0);
    rms_norm_16_div_cmp_z : IN STD_LOGIC_VECTOR (71 DOWNTO 0);
    attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_pff : OUT STD_LOGIC;
    attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_pff : OUT STD_LOGIC;
    attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_pff : OUT STD_LOGIC;
    attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_pff : OUT STD_LOGIC;
    attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_pff : OUT STD_LOGIC
  );
END dut_core;

ARCHITECTURE v1 OF dut_core IS
  -- Interconnect Declarations
  SIGNAL core_wen1 : STD_LOGIC;
  SIGNAL strm_in_rsci_wen_comp : STD_LOGIC;
  SIGNAL strm_in_rsci_idat_mxwt : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL strm_out_rsci_wen_comp : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 : STD_LOGIC;
  SIGNAL SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z : STD_LOGIC_VECTOR (55 DOWNTO
      0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z
      : STD_LOGIC_VECTOR (71 DOWNTO 0);
  SIGNAL rms_norm_16_div_cmp_z_oreg : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_71_48
      : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL strm_out_rsci_idat_31_18 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL fsm_output : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_2_2_acc_1_tmp : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CM_LOOP_3_acc_tmp : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_acc_6_tmp : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL CACHE_UPDATE_LOOP_1_and_tmp : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL for_for_and_tmp : STD_LOGIC;
  SIGNAL or_dcpl_4 : STD_LOGIC;
  SIGNAL and_dcpl : STD_LOGIC;
  SIGNAL and_dcpl_1 : STD_LOGIC;
  SIGNAL or_tmp_11 : STD_LOGIC;
  SIGNAL or_tmp_48 : STD_LOGIC;
  SIGNAL or_dcpl_45 : STD_LOGIC;
  SIGNAL or_dcpl_47 : STD_LOGIC;
  SIGNAL or_dcpl_54 : STD_LOGIC;
  SIGNAL or_dcpl_60 : STD_LOGIC;
  SIGNAL or_dcpl_68 : STD_LOGIC;
  SIGNAL or_dcpl_79 : STD_LOGIC;
  SIGNAL or_dcpl_96 : STD_LOGIC;
  SIGNAL or_tmp_104 : STD_LOGIC;
  SIGNAL mux_tmp_87 : STD_LOGIC;
  SIGNAL mux_tmp_91 : STD_LOGIC;
  SIGNAL nor_tmp_28 : STD_LOGIC;
  SIGNAL mux_tmp_121 : STD_LOGIC;
  SIGNAL and_dcpl_26 : STD_LOGIC;
  SIGNAL and_dcpl_45 : STD_LOGIC;
  SIGNAL nor_tmp_99 : STD_LOGIC;
  SIGNAL and_dcpl_57 : STD_LOGIC;
  SIGNAL and_dcpl_61 : STD_LOGIC;
  SIGNAL and_dcpl_65 : STD_LOGIC;
  SIGNAL or_dcpl_332 : STD_LOGIC;
  SIGNAL or_dcpl_337 : STD_LOGIC;
  SIGNAL or_dcpl_342 : STD_LOGIC;
  SIGNAL or_dcpl_351 : STD_LOGIC;
  SIGNAL or_dcpl_377 : STD_LOGIC;
  SIGNAL or_tmp_330 : STD_LOGIC;
  SIGNAL nor_tmp_117 : STD_LOGIC;
  SIGNAL mux_tmp_363 : STD_LOGIC;
  SIGNAL not_tmp_253 : STD_LOGIC;
  SIGNAL or_dcpl_508 : STD_LOGIC;
  SIGNAL or_dcpl_512 : STD_LOGIC;
  SIGNAL or_dcpl_584 : STD_LOGIC;
  SIGNAL or_tmp_464 : STD_LOGIC;
  SIGNAL or_dcpl_672 : STD_LOGIC;
  SIGNAL or_tmp_507 : STD_LOGIC;
  SIGNAL mux_tmp_604 : STD_LOGIC;
  SIGNAL or_tmp_611 : STD_LOGIC;
  SIGNAL or_dcpl_770 : STD_LOGIC;
  SIGNAL or_dcpl_774 : STD_LOGIC;
  SIGNAL or_dcpl_791 : STD_LOGIC;
  SIGNAL or_dcpl_794 : STD_LOGIC;
  SIGNAL and_dcpl_148 : STD_LOGIC;
  SIGNAL or_tmp_682 : STD_LOGIC;
  SIGNAL or_dcpl_959 : STD_LOGIC;
  SIGNAL or_dcpl_961 : STD_LOGIC;
  SIGNAL and_dcpl_181 : STD_LOGIC;
  SIGNAL and_dcpl_182 : STD_LOGIC;
  SIGNAL and_dcpl_185 : STD_LOGIC;
  SIGNAL and_dcpl_186 : STD_LOGIC;
  SIGNAL and_dcpl_187 : STD_LOGIC;
  SIGNAL and_dcpl_189 : STD_LOGIC;
  SIGNAL and_dcpl_190 : STD_LOGIC;
  SIGNAL and_dcpl_191 : STD_LOGIC;
  SIGNAL and_dcpl_192 : STD_LOGIC;
  SIGNAL and_dcpl_193 : STD_LOGIC;
  SIGNAL and_dcpl_194 : STD_LOGIC;
  SIGNAL and_dcpl_197 : STD_LOGIC;
  SIGNAL and_dcpl_198 : STD_LOGIC;
  SIGNAL and_dcpl_199 : STD_LOGIC;
  SIGNAL and_dcpl_200 : STD_LOGIC;
  SIGNAL and_dcpl_201 : STD_LOGIC;
  SIGNAL and_dcpl_202 : STD_LOGIC;
  SIGNAL and_dcpl_203 : STD_LOGIC;
  SIGNAL and_dcpl_204 : STD_LOGIC;
  SIGNAL or_dcpl_980 : STD_LOGIC;
  SIGNAL or_dcpl_983 : STD_LOGIC;
  SIGNAL or_dcpl_985 : STD_LOGIC;
  SIGNAL or_dcpl_987 : STD_LOGIC;
  SIGNAL or_dcpl_988 : STD_LOGIC;
  SIGNAL or_dcpl_989 : STD_LOGIC;
  SIGNAL or_dcpl_990 : STD_LOGIC;
  SIGNAL or_dcpl_991 : STD_LOGIC;
  SIGNAL or_dcpl_993 : STD_LOGIC;
  SIGNAL or_dcpl_995 : STD_LOGIC;
  SIGNAL or_dcpl_996 : STD_LOGIC;
  SIGNAL or_dcpl_997 : STD_LOGIC;
  SIGNAL or_dcpl_998 : STD_LOGIC;
  SIGNAL or_dcpl_999 : STD_LOGIC;
  SIGNAL or_dcpl_1000 : STD_LOGIC;
  SIGNAL and_dcpl_205 : STD_LOGIC;
  SIGNAL and_dcpl_206 : STD_LOGIC;
  SIGNAL and_dcpl_207 : STD_LOGIC;
  SIGNAL or_dcpl_1001 : STD_LOGIC;
  SIGNAL or_dcpl_1002 : STD_LOGIC;
  SIGNAL or_dcpl_1003 : STD_LOGIC;
  SIGNAL or_dcpl_1004 : STD_LOGIC;
  SIGNAL or_dcpl_1005 : STD_LOGIC;
  SIGNAL or_dcpl_1006 : STD_LOGIC;
  SIGNAL or_dcpl_1007 : STD_LOGIC;
  SIGNAL or_dcpl_1008 : STD_LOGIC;
  SIGNAL or_dcpl_1009 : STD_LOGIC;
  SIGNAL or_dcpl_1010 : STD_LOGIC;
  SIGNAL or_dcpl_1011 : STD_LOGIC;
  SIGNAL or_dcpl_1012 : STD_LOGIC;
  SIGNAL or_dcpl_1013 : STD_LOGIC;
  SIGNAL or_dcpl_1014 : STD_LOGIC;
  SIGNAL or_dcpl_1015 : STD_LOGIC;
  SIGNAL or_dcpl_1016 : STD_LOGIC;
  SIGNAL or_dcpl_1017 : STD_LOGIC;
  SIGNAL or_dcpl_1018 : STD_LOGIC;
  SIGNAL or_dcpl_1019 : STD_LOGIC;
  SIGNAL and_dcpl_209 : STD_LOGIC;
  SIGNAL and_dcpl_211 : STD_LOGIC;
  SIGNAL and_dcpl_212 : STD_LOGIC;
  SIGNAL and_dcpl_213 : STD_LOGIC;
  SIGNAL nor_tmp_261 : STD_LOGIC;
  SIGNAL and_dcpl_215 : STD_LOGIC;
  SIGNAL and_dcpl_216 : STD_LOGIC;
  SIGNAL mux_tmp_787 : STD_LOGIC;
  SIGNAL mux_tmp_788 : STD_LOGIC;
  SIGNAL and_dcpl_220 : STD_LOGIC;
  SIGNAL and_dcpl_221 : STD_LOGIC;
  SIGNAL and_dcpl_222 : STD_LOGIC;
  SIGNAL or_dcpl_1020 : STD_LOGIC;
  SIGNAL or_dcpl_1021 : STD_LOGIC;
  SIGNAL or_dcpl_1022 : STD_LOGIC;
  SIGNAL or_dcpl_1023 : STD_LOGIC;
  SIGNAL or_dcpl_1024 : STD_LOGIC;
  SIGNAL and_dcpl_226 : STD_LOGIC;
  SIGNAL or_tmp_704 : STD_LOGIC;
  SIGNAL or_tmp_708 : STD_LOGIC;
  SIGNAL and_dcpl_231 : STD_LOGIC;
  SIGNAL or_dcpl_1025 : STD_LOGIC;
  SIGNAL and_dcpl_237 : STD_LOGIC;
  SIGNAL and_dcpl_239 : STD_LOGIC;
  SIGNAL and_dcpl_240 : STD_LOGIC;
  SIGNAL or_dcpl_1026 : STD_LOGIC;
  SIGNAL or_dcpl_1027 : STD_LOGIC;
  SIGNAL or_dcpl_1028 : STD_LOGIC;
  SIGNAL or_dcpl_1029 : STD_LOGIC;
  SIGNAL or_dcpl_1030 : STD_LOGIC;
  SIGNAL or_dcpl_1031 : STD_LOGIC;
  SIGNAL or_dcpl_1032 : STD_LOGIC;
  SIGNAL or_dcpl_1033 : STD_LOGIC;
  SIGNAL or_dcpl_1034 : STD_LOGIC;
  SIGNAL or_dcpl_1035 : STD_LOGIC;
  SIGNAL or_dcpl_1036 : STD_LOGIC;
  SIGNAL or_dcpl_1037 : STD_LOGIC;
  SIGNAL or_dcpl_1038 : STD_LOGIC;
  SIGNAL or_dcpl_1039 : STD_LOGIC;
  SIGNAL or_dcpl_1040 : STD_LOGIC;
  SIGNAL or_dcpl_1041 : STD_LOGIC;
  SIGNAL or_dcpl_1042 : STD_LOGIC;
  SIGNAL or_dcpl_1043 : STD_LOGIC;
  SIGNAL or_dcpl_1044 : STD_LOGIC;
  SIGNAL or_dcpl_1045 : STD_LOGIC;
  SIGNAL or_dcpl_1046 : STD_LOGIC;
  SIGNAL and_dcpl_241 : STD_LOGIC;
  SIGNAL and_dcpl_242 : STD_LOGIC;
  SIGNAL and_dcpl_243 : STD_LOGIC;
  SIGNAL and_dcpl_248 : STD_LOGIC;
  SIGNAL and_dcpl_252 : STD_LOGIC;
  SIGNAL and_dcpl_255 : STD_LOGIC;
  SIGNAL and_dcpl_256 : STD_LOGIC;
  SIGNAL and_dcpl_257 : STD_LOGIC;
  SIGNAL and_dcpl_258 : STD_LOGIC;
  SIGNAL and_dcpl_259 : STD_LOGIC;
  SIGNAL or_tmp_728 : STD_LOGIC;
  SIGNAL and_dcpl_260 : STD_LOGIC;
  SIGNAL mux_tmp_824 : STD_LOGIC;
  SIGNAL or_dcpl_1048 : STD_LOGIC;
  SIGNAL and_dcpl_261 : STD_LOGIC;
  SIGNAL and_dcpl_263 : STD_LOGIC;
  SIGNAL and_dcpl_264 : STD_LOGIC;
  SIGNAL and_dcpl_265 : STD_LOGIC;
  SIGNAL or_dcpl_1050 : STD_LOGIC;
  SIGNAL and_dcpl_268 : STD_LOGIC;
  SIGNAL and_dcpl_270 : STD_LOGIC;
  SIGNAL mux_tmp_834 : STD_LOGIC;
  SIGNAL mux_tmp_836 : STD_LOGIC;
  SIGNAL and_dcpl_272 : STD_LOGIC;
  SIGNAL and_dcpl_275 : STD_LOGIC;
  SIGNAL and_dcpl_276 : STD_LOGIC;
  SIGNAL nor_tmp_282 : STD_LOGIC;
  SIGNAL and_dcpl_278 : STD_LOGIC;
  SIGNAL and_dcpl_279 : STD_LOGIC;
  SIGNAL or_tmp_742 : STD_LOGIC;
  SIGNAL mux_tmp_839 : STD_LOGIC;
  SIGNAL mux_tmp_841 : STD_LOGIC;
  SIGNAL nor_tmp_285 : STD_LOGIC;
  SIGNAL and_dcpl_289 : STD_LOGIC;
  SIGNAL and_dcpl_290 : STD_LOGIC;
  SIGNAL and_dcpl_291 : STD_LOGIC;
  SIGNAL and_dcpl_292 : STD_LOGIC;
  SIGNAL and_dcpl_293 : STD_LOGIC;
  SIGNAL and_dcpl_294 : STD_LOGIC;
  SIGNAL and_dcpl_295 : STD_LOGIC;
  SIGNAL or_tmp_755 : STD_LOGIC;
  SIGNAL and_dcpl_298 : STD_LOGIC;
  SIGNAL and_dcpl_302 : STD_LOGIC;
  SIGNAL or_tmp_757 : STD_LOGIC;
  SIGNAL or_tmp_762 : STD_LOGIC;
  SIGNAL mux_tmp_857 : STD_LOGIC;
  SIGNAL and_dcpl_304 : STD_LOGIC;
  SIGNAL nor_tmp_289 : STD_LOGIC;
  SIGNAL and_dcpl_306 : STD_LOGIC;
  SIGNAL and_dcpl_307 : STD_LOGIC;
  SIGNAL and_dcpl_308 : STD_LOGIC;
  SIGNAL nor_tmp_291 : STD_LOGIC;
  SIGNAL or_tmp_767 : STD_LOGIC;
  SIGNAL and_dcpl_310 : STD_LOGIC;
  SIGNAL and_dcpl_312 : STD_LOGIC;
  SIGNAL and_dcpl_313 : STD_LOGIC;
  SIGNAL and_dcpl_315 : STD_LOGIC;
  SIGNAL and_dcpl_316 : STD_LOGIC;
  SIGNAL and_dcpl_318 : STD_LOGIC;
  SIGNAL and_dcpl_319 : STD_LOGIC;
  SIGNAL and_dcpl_321 : STD_LOGIC;
  SIGNAL and_dcpl_322 : STD_LOGIC;
  SIGNAL and_dcpl_327 : STD_LOGIC;
  SIGNAL and_dcpl_328 : STD_LOGIC;
  SIGNAL and_dcpl_334 : STD_LOGIC;
  SIGNAL and_dcpl_335 : STD_LOGIC;
  SIGNAL and_dcpl_336 : STD_LOGIC;
  SIGNAL and_dcpl_338 : STD_LOGIC;
  SIGNAL and_dcpl_339 : STD_LOGIC;
  SIGNAL and_dcpl_341 : STD_LOGIC;
  SIGNAL and_dcpl_342 : STD_LOGIC;
  SIGNAL nor_tmp_307 : STD_LOGIC;
  SIGNAL and_dcpl_344 : STD_LOGIC;
  SIGNAL and_dcpl_346 : STD_LOGIC;
  SIGNAL or_tmp_798 : STD_LOGIC;
  SIGNAL and_dcpl_348 : STD_LOGIC;
  SIGNAL and_dcpl_349 : STD_LOGIC;
  SIGNAL and_dcpl_350 : STD_LOGIC;
  SIGNAL and_dcpl_351 : STD_LOGIC;
  SIGNAL and_dcpl_352 : STD_LOGIC;
  SIGNAL and_dcpl_353 : STD_LOGIC;
  SIGNAL and_dcpl_354 : STD_LOGIC;
  SIGNAL and_dcpl_355 : STD_LOGIC;
  SIGNAL and_dcpl_357 : STD_LOGIC;
  SIGNAL and_dcpl_360 : STD_LOGIC;
  SIGNAL or_dcpl_1063 : STD_LOGIC;
  SIGNAL and_dcpl_362 : STD_LOGIC;
  SIGNAL and_dcpl_363 : STD_LOGIC;
  SIGNAL and_dcpl_364 : STD_LOGIC;
  SIGNAL and_dcpl_374 : STD_LOGIC;
  SIGNAL or_tmp_805 : STD_LOGIC;
  SIGNAL mux_tmp_906 : STD_LOGIC;
  SIGNAL or_tmp_808 : STD_LOGIC;
  SIGNAL mux_tmp_908 : STD_LOGIC;
  SIGNAL mux_tmp_910 : STD_LOGIC;
  SIGNAL or_tmp_812 : STD_LOGIC;
  SIGNAL mux_tmp_915 : STD_LOGIC;
  SIGNAL or_tmp_813 : STD_LOGIC;
  SIGNAL mux_tmp_916 : STD_LOGIC;
  SIGNAL mux_tmp_919 : STD_LOGIC;
  SIGNAL or_tmp_814 : STD_LOGIC;
  SIGNAL mux_tmp_922 : STD_LOGIC;
  SIGNAL mux_tmp_927 : STD_LOGIC;
  SIGNAL mux_tmp_936 : STD_LOGIC;
  SIGNAL mux_tmp_937 : STD_LOGIC;
  SIGNAL and_dcpl_376 : STD_LOGIC;
  SIGNAL and_dcpl_377 : STD_LOGIC;
  SIGNAL and_dcpl_381 : STD_LOGIC;
  SIGNAL and_dcpl_382 : STD_LOGIC;
  SIGNAL or_tmp_833 : STD_LOGIC;
  SIGNAL mux_tmp_960 : STD_LOGIC;
  SIGNAL mux_tmp_967 : STD_LOGIC;
  SIGNAL mux_tmp_968 : STD_LOGIC;
  SIGNAL and_dcpl_383 : STD_LOGIC;
  SIGNAL mux_tmp_975 : STD_LOGIC;
  SIGNAL and_dcpl_385 : STD_LOGIC;
  SIGNAL and_dcpl_386 : STD_LOGIC;
  SIGNAL and_dcpl_388 : STD_LOGIC;
  SIGNAL or_tmp_861 : STD_LOGIC;
  SIGNAL and_dcpl_390 : STD_LOGIC;
  SIGNAL or_tmp_878 : STD_LOGIC;
  SIGNAL and_dcpl_410 : STD_LOGIC;
  SIGNAL and_dcpl_413 : STD_LOGIC;
  SIGNAL nor_tmp_329 : STD_LOGIC;
  SIGNAL mux_tmp_1027 : STD_LOGIC;
  SIGNAL and_dcpl_414 : STD_LOGIC;
  SIGNAL and_dcpl_415 : STD_LOGIC;
  SIGNAL or_tmp_913 : STD_LOGIC;
  SIGNAL or_tmp_914 : STD_LOGIC;
  SIGNAL and_dcpl_417 : STD_LOGIC;
  SIGNAL and_dcpl_420 : STD_LOGIC;
  SIGNAL and_dcpl_421 : STD_LOGIC;
  SIGNAL and_dcpl_422 : STD_LOGIC;
  SIGNAL or_dcpl_1067 : STD_LOGIC;
  SIGNAL and_dcpl_425 : STD_LOGIC;
  SIGNAL or_tmp_922 : STD_LOGIC;
  SIGNAL or_tmp_923 : STD_LOGIC;
  SIGNAL mux_tmp_1044 : STD_LOGIC;
  SIGNAL or_tmp_930 : STD_LOGIC;
  SIGNAL mux_tmp_1051 : STD_LOGIC;
  SIGNAL mux_tmp_1052 : STD_LOGIC;
  SIGNAL or_tmp_931 : STD_LOGIC;
  SIGNAL or_dcpl_1068 : STD_LOGIC;
  SIGNAL and_dcpl_432 : STD_LOGIC;
  SIGNAL and_dcpl_433 : STD_LOGIC;
  SIGNAL or_dcpl_1070 : STD_LOGIC;
  SIGNAL or_dcpl_1071 : STD_LOGIC;
  SIGNAL and_dcpl_438 : STD_LOGIC;
  SIGNAL and_dcpl_439 : STD_LOGIC;
  SIGNAL or_tmp_938 : STD_LOGIC;
  SIGNAL not_tmp_549 : STD_LOGIC;
  SIGNAL and_dcpl_442 : STD_LOGIC;
  SIGNAL and_dcpl_448 : STD_LOGIC;
  SIGNAL and_dcpl_449 : STD_LOGIC;
  SIGNAL and_dcpl_452 : STD_LOGIC;
  SIGNAL and_dcpl_453 : STD_LOGIC;
  SIGNAL or_dcpl_1073 : STD_LOGIC;
  SIGNAL and_dcpl_458 : STD_LOGIC;
  SIGNAL or_dcpl_1076 : STD_LOGIC;
  SIGNAL and_dcpl_461 : STD_LOGIC;
  SIGNAL and_dcpl_462 : STD_LOGIC;
  SIGNAL or_dcpl_1077 : STD_LOGIC;
  SIGNAL or_dcpl_1079 : STD_LOGIC;
  SIGNAL and_dcpl_467 : STD_LOGIC;
  SIGNAL and_dcpl_468 : STD_LOGIC;
  SIGNAL or_dcpl_1081 : STD_LOGIC;
  SIGNAL and_dcpl_471 : STD_LOGIC;
  SIGNAL or_dcpl_1083 : STD_LOGIC;
  SIGNAL and_dcpl_477 : STD_LOGIC;
  SIGNAL and_dcpl_478 : STD_LOGIC;
  SIGNAL or_tmp_992 : STD_LOGIC;
  SIGNAL mux_tmp_1113 : STD_LOGIC;
  SIGNAL or_tmp_993 : STD_LOGIC;
  SIGNAL and_dcpl_480 : STD_LOGIC;
  SIGNAL or_dcpl_1084 : STD_LOGIC;
  SIGNAL and_dcpl_486 : STD_LOGIC;
  SIGNAL or_dcpl_1085 : STD_LOGIC;
  SIGNAL or_dcpl_1086 : STD_LOGIC;
  SIGNAL or_dcpl_1087 : STD_LOGIC;
  SIGNAL or_dcpl_1088 : STD_LOGIC;
  SIGNAL or_dcpl_1089 : STD_LOGIC;
  SIGNAL mux_tmp_1120 : STD_LOGIC;
  SIGNAL and_dcpl_511 : STD_LOGIC;
  SIGNAL and_dcpl_512 : STD_LOGIC;
  SIGNAL and_dcpl_513 : STD_LOGIC;
  SIGNAL or_dcpl_1090 : STD_LOGIC;
  SIGNAL and_dcpl_524 : STD_LOGIC;
  SIGNAL mux_tmp_1163 : STD_LOGIC;
  SIGNAL and_dcpl_525 : STD_LOGIC;
  SIGNAL and_dcpl_528 : STD_LOGIC;
  SIGNAL or_dcpl_1091 : STD_LOGIC;
  SIGNAL or_dcpl_1092 : STD_LOGIC;
  SIGNAL mux_tmp_1178 : STD_LOGIC;
  SIGNAL mux_tmp_1179 : STD_LOGIC;
  SIGNAL mux_tmp_1183 : STD_LOGIC;
  SIGNAL mux_tmp_1185 : STD_LOGIC;
  SIGNAL mux_tmp_1187 : STD_LOGIC;
  SIGNAL or_tmp_1035 : STD_LOGIC;
  SIGNAL and_dcpl_539 : STD_LOGIC;
  SIGNAL or_tmp_1051 : STD_LOGIC;
  SIGNAL mux_tmp_1218 : STD_LOGIC;
  SIGNAL mux_tmp_1219 : STD_LOGIC;
  SIGNAL mux_tmp_1229 : STD_LOGIC;
  SIGNAL mux_tmp_1237 : STD_LOGIC;
  SIGNAL mux_tmp_1238 : STD_LOGIC;
  SIGNAL or_tmp_1066 : STD_LOGIC;
  SIGNAL mux_tmp_1240 : STD_LOGIC;
  SIGNAL mux_tmp_1245 : STD_LOGIC;
  SIGNAL mux_tmp_1250 : STD_LOGIC;
  SIGNAL and_dcpl_548 : STD_LOGIC;
  SIGNAL and_dcpl_549 : STD_LOGIC;
  SIGNAL and_dcpl_550 : STD_LOGIC;
  SIGNAL and_dcpl_551 : STD_LOGIC;
  SIGNAL and_dcpl_552 : STD_LOGIC;
  SIGNAL and_dcpl_553 : STD_LOGIC;
  SIGNAL and_dcpl_554 : STD_LOGIC;
  SIGNAL and_dcpl_557 : STD_LOGIC;
  SIGNAL mux_tmp_1281 : STD_LOGIC;
  SIGNAL and_dcpl_564 : STD_LOGIC;
  SIGNAL and_dcpl_576 : STD_LOGIC;
  SIGNAL and_dcpl_577 : STD_LOGIC;
  SIGNAL and_dcpl_581 : STD_LOGIC;
  SIGNAL or_tmp_1128 : STD_LOGIC;
  SIGNAL and_dcpl_583 : STD_LOGIC;
  SIGNAL or_tmp_1132 : STD_LOGIC;
  SIGNAL or_dcpl_1104 : STD_LOGIC;
  SIGNAL and_dcpl_585 : STD_LOGIC;
  SIGNAL and_dcpl_586 : STD_LOGIC;
  SIGNAL and_dcpl_587 : STD_LOGIC;
  SIGNAL and_dcpl_588 : STD_LOGIC;
  SIGNAL and_dcpl_591 : STD_LOGIC;
  SIGNAL and_dcpl_592 : STD_LOGIC;
  SIGNAL and_dcpl_595 : STD_LOGIC;
  SIGNAL and_dcpl_598 : STD_LOGIC;
  SIGNAL and_dcpl_601 : STD_LOGIC;
  SIGNAL and_dcpl_604 : STD_LOGIC;
  SIGNAL and_dcpl_607 : STD_LOGIC;
  SIGNAL and_dcpl_610 : STD_LOGIC;
  SIGNAL and_dcpl_613 : STD_LOGIC;
  SIGNAL and_dcpl_616 : STD_LOGIC;
  SIGNAL and_dcpl_618 : STD_LOGIC;
  SIGNAL and_dcpl_619 : STD_LOGIC;
  SIGNAL or_tmp_1203 : STD_LOGIC;
  SIGNAL and_dcpl_620 : STD_LOGIC;
  SIGNAL mux_tmp_1421 : STD_LOGIC;
  SIGNAL or_tmp_1218 : STD_LOGIC;
  SIGNAL not_tmp_650 : STD_LOGIC;
  SIGNAL and_dcpl_622 : STD_LOGIC;
  SIGNAL and_dcpl_625 : STD_LOGIC;
  SIGNAL or_tmp_1221 : STD_LOGIC;
  SIGNAL mux_tmp_1426 : STD_LOGIC;
  SIGNAL and_dcpl_626 : STD_LOGIC;
  SIGNAL and_dcpl_628 : STD_LOGIC;
  SIGNAL and_dcpl_629 : STD_LOGIC;
  SIGNAL mux_tmp_1440 : STD_LOGIC;
  SIGNAL and_dcpl_635 : STD_LOGIC;
  SIGNAL and_tmp_42 : STD_LOGIC;
  SIGNAL mux_tmp_1451 : STD_LOGIC;
  SIGNAL and_dcpl_641 : STD_LOGIC;
  SIGNAL and_dcpl_642 : STD_LOGIC;
  SIGNAL or_dcpl_1108 : STD_LOGIC;
  SIGNAL mux_tmp_1489 : STD_LOGIC;
  SIGNAL or_dcpl_1109 : STD_LOGIC;
  SIGNAL or_dcpl_1114 : STD_LOGIC;
  SIGNAL and_dcpl_650 : STD_LOGIC;
  SIGNAL and_dcpl_651 : STD_LOGIC;
  SIGNAL or_dcpl_1116 : STD_LOGIC;
  SIGNAL and_dcpl_656 : STD_LOGIC;
  SIGNAL or_dcpl_1118 : STD_LOGIC;
  SIGNAL or_dcpl_1119 : STD_LOGIC;
  SIGNAL or_dcpl_1120 : STD_LOGIC;
  SIGNAL or_dcpl_1121 : STD_LOGIC;
  SIGNAL or_dcpl_1122 : STD_LOGIC;
  SIGNAL or_dcpl_1123 : STD_LOGIC;
  SIGNAL or_dcpl_1125 : STD_LOGIC;
  SIGNAL or_dcpl_1126 : STD_LOGIC;
  SIGNAL or_dcpl_1127 : STD_LOGIC;
  SIGNAL or_dcpl_1128 : STD_LOGIC;
  SIGNAL or_dcpl_1130 : STD_LOGIC;
  SIGNAL or_dcpl_1131 : STD_LOGIC;
  SIGNAL or_dcpl_1132 : STD_LOGIC;
  SIGNAL or_dcpl_1133 : STD_LOGIC;
  SIGNAL or_tmp_1291 : STD_LOGIC;
  SIGNAL or_tmp_1296 : STD_LOGIC;
  SIGNAL and_dcpl_718 : STD_LOGIC;
  SIGNAL or_tmp_1316 : STD_LOGIC;
  SIGNAL mux_tmp_1519 : STD_LOGIC;
  SIGNAL or_tmp_1320 : STD_LOGIC;
  SIGNAL and_dcpl_721 : STD_LOGIC;
  SIGNAL not_tmp_699 : STD_LOGIC;
  SIGNAL and_dcpl_725 : STD_LOGIC;
  SIGNAL and_dcpl_726 : STD_LOGIC;
  SIGNAL or_dcpl_1134 : STD_LOGIC;
  SIGNAL or_dcpl_1137 : STD_LOGIC;
  SIGNAL or_dcpl_1138 : STD_LOGIC;
  SIGNAL or_dcpl_1140 : STD_LOGIC;
  SIGNAL or_dcpl_1141 : STD_LOGIC;
  SIGNAL and_dcpl_727 : STD_LOGIC;
  SIGNAL and_dcpl_728 : STD_LOGIC;
  SIGNAL and_dcpl_729 : STD_LOGIC;
  SIGNAL and_dcpl_730 : STD_LOGIC;
  SIGNAL and_dcpl_731 : STD_LOGIC;
  SIGNAL and_dcpl_732 : STD_LOGIC;
  SIGNAL mux_tmp_1548 : STD_LOGIC;
  SIGNAL mux_tmp_1549 : STD_LOGIC;
  SIGNAL nand_tmp_66 : STD_LOGIC;
  SIGNAL and_dcpl_735 : STD_LOGIC;
  SIGNAL and_dcpl_736 : STD_LOGIC;
  SIGNAL and_dcpl_739 : STD_LOGIC;
  SIGNAL and_dcpl_740 : STD_LOGIC;
  SIGNAL and_dcpl_743 : STD_LOGIC;
  SIGNAL and_dcpl_745 : STD_LOGIC;
  SIGNAL and_dcpl_747 : STD_LOGIC;
  SIGNAL and_dcpl_748 : STD_LOGIC;
  SIGNAL mux_tmp_1562 : STD_LOGIC;
  SIGNAL and_dcpl_751 : STD_LOGIC;
  SIGNAL and_dcpl_753 : STD_LOGIC;
  SIGNAL and_dcpl_754 : STD_LOGIC;
  SIGNAL and_dcpl_758 : STD_LOGIC;
  SIGNAL and_dcpl_760 : STD_LOGIC;
  SIGNAL and_dcpl_764 : STD_LOGIC;
  SIGNAL and_dcpl_768 : STD_LOGIC;
  SIGNAL and_dcpl_772 : STD_LOGIC;
  SIGNAL and_dcpl_776 : STD_LOGIC;
  SIGNAL and_dcpl_780 : STD_LOGIC;
  SIGNAL and_dcpl_784 : STD_LOGIC;
  SIGNAL and_dcpl_788 : STD_LOGIC;
  SIGNAL and_dcpl_792 : STD_LOGIC;
  SIGNAL and_dcpl_796 : STD_LOGIC;
  SIGNAL and_dcpl_800 : STD_LOGIC;
  SIGNAL and_dcpl_804 : STD_LOGIC;
  SIGNAL and_dcpl_810 : STD_LOGIC;
  SIGNAL and_dcpl_812 : STD_LOGIC;
  SIGNAL and_dcpl_813 : STD_LOGIC;
  SIGNAL and_dcpl_814 : STD_LOGIC;
  SIGNAL mux_tmp_1578 : STD_LOGIC;
  SIGNAL and_dcpl_817 : STD_LOGIC;
  SIGNAL and_dcpl_818 : STD_LOGIC;
  SIGNAL and_dcpl_819 : STD_LOGIC;
  SIGNAL and_dcpl_820 : STD_LOGIC;
  SIGNAL and_dcpl_821 : STD_LOGIC;
  SIGNAL or_tmp_1354 : STD_LOGIC;
  SIGNAL and_dcpl_825 : STD_LOGIC;
  SIGNAL and_dcpl_826 : STD_LOGIC;
  SIGNAL and_dcpl_827 : STD_LOGIC;
  SIGNAL and_dcpl_830 : STD_LOGIC;
  SIGNAL and_dcpl_831 : STD_LOGIC;
  SIGNAL and_dcpl_832 : STD_LOGIC;
  SIGNAL and_dcpl_835 : STD_LOGIC;
  SIGNAL and_dcpl_836 : STD_LOGIC;
  SIGNAL and_dcpl_837 : STD_LOGIC;
  SIGNAL and_dcpl_840 : STD_LOGIC;
  SIGNAL and_dcpl_841 : STD_LOGIC;
  SIGNAL and_dcpl_842 : STD_LOGIC;
  SIGNAL and_dcpl_843 : STD_LOGIC;
  SIGNAL and_dcpl_847 : STD_LOGIC;
  SIGNAL and_dcpl_850 : STD_LOGIC;
  SIGNAL and_dcpl_851 : STD_LOGIC;
  SIGNAL and_dcpl_854 : STD_LOGIC;
  SIGNAL and_dcpl_855 : STD_LOGIC;
  SIGNAL and_dcpl_856 : STD_LOGIC;
  SIGNAL and_dcpl_859 : STD_LOGIC;
  SIGNAL and_dcpl_860 : STD_LOGIC;
  SIGNAL and_dcpl_863 : STD_LOGIC;
  SIGNAL and_dcpl_864 : STD_LOGIC;
  SIGNAL and_dcpl_867 : STD_LOGIC;
  SIGNAL and_dcpl_868 : STD_LOGIC;
  SIGNAL and_dcpl_871 : STD_LOGIC;
  SIGNAL and_dcpl_872 : STD_LOGIC;
  SIGNAL and_dcpl_875 : STD_LOGIC;
  SIGNAL and_dcpl_876 : STD_LOGIC;
  SIGNAL and_dcpl_879 : STD_LOGIC;
  SIGNAL and_dcpl_880 : STD_LOGIC;
  SIGNAL and_dcpl_885 : STD_LOGIC;
  SIGNAL or_tmp_1392 : STD_LOGIC;
  SIGNAL and_dcpl_888 : STD_LOGIC;
  SIGNAL and_dcpl_959 : STD_LOGIC;
  SIGNAL mux_tmp_1943 : STD_LOGIC;
  SIGNAL mux_tmp_1945 : STD_LOGIC;
  SIGNAL and_dcpl_983 : STD_LOGIC;
  SIGNAL and_dcpl_987 : STD_LOGIC;
  SIGNAL and_dcpl_989 : STD_LOGIC;
  SIGNAL and_dcpl_999 : STD_LOGIC;
  SIGNAL and_dcpl_1000 : STD_LOGIC;
  SIGNAL mux_tmp_1990 : STD_LOGIC;
  SIGNAL mux_tmp_1993 : STD_LOGIC;
  SIGNAL and_dcpl_1003 : STD_LOGIC;
  SIGNAL or_dcpl_1145 : STD_LOGIC;
  SIGNAL mux_tmp_2013 : STD_LOGIC;
  SIGNAL mux_tmp_2015 : STD_LOGIC;
  SIGNAL or_dcpl_1146 : STD_LOGIC;
  SIGNAL mux_tmp_2034 : STD_LOGIC;
  SIGNAL and_dcpl_1011 : STD_LOGIC;
  SIGNAL and_dcpl_1033 : STD_LOGIC;
  SIGNAL and_dcpl_1034 : STD_LOGIC;
  SIGNAL mux_tmp_2067 : STD_LOGIC;
  SIGNAL and_dcpl_1055 : STD_LOGIC;
  SIGNAL and_dcpl_1061 : STD_LOGIC;
  SIGNAL or_tmp_1632 : STD_LOGIC;
  SIGNAL not_tmp_874 : STD_LOGIC;
  SIGNAL or_tmp_1643 : STD_LOGIC;
  SIGNAL or_dcpl_1152 : STD_LOGIC;
  SIGNAL or_dcpl_1155 : STD_LOGIC;
  SIGNAL or_dcpl_1156 : STD_LOGIC;
  SIGNAL or_dcpl_1158 : STD_LOGIC;
  SIGNAL or_dcpl_1159 : STD_LOGIC;
  SIGNAL or_dcpl_1160 : STD_LOGIC;
  SIGNAL or_dcpl_1161 : STD_LOGIC;
  SIGNAL or_dcpl_1162 : STD_LOGIC;
  SIGNAL or_dcpl_1163 : STD_LOGIC;
  SIGNAL or_dcpl_1164 : STD_LOGIC;
  SIGNAL or_dcpl_1165 : STD_LOGIC;
  SIGNAL or_dcpl_1166 : STD_LOGIC;
  SIGNAL or_dcpl_1167 : STD_LOGIC;
  SIGNAL or_dcpl_1168 : STD_LOGIC;
  SIGNAL or_dcpl_1169 : STD_LOGIC;
  SIGNAL or_dcpl_1170 : STD_LOGIC;
  SIGNAL and_dcpl_1073 : STD_LOGIC;
  SIGNAL and_dcpl_1082 : STD_LOGIC;
  SIGNAL and_dcpl_1084 : STD_LOGIC;
  SIGNAL and_dcpl_1088 : STD_LOGIC;
  SIGNAL and_dcpl_1091 : STD_LOGIC;
  SIGNAL and_dcpl_1094 : STD_LOGIC;
  SIGNAL and_dcpl_1097 : STD_LOGIC;
  SIGNAL and_dcpl_1100 : STD_LOGIC;
  SIGNAL and_dcpl_1103 : STD_LOGIC;
  SIGNAL and_dcpl_1106 : STD_LOGIC;
  SIGNAL and_dcpl_1109 : STD_LOGIC;
  SIGNAL and_dcpl_1112 : STD_LOGIC;
  SIGNAL and_dcpl_1115 : STD_LOGIC;
  SIGNAL and_dcpl_1118 : STD_LOGIC;
  SIGNAL and_dcpl_1121 : STD_LOGIC;
  SIGNAL and_dcpl_1124 : STD_LOGIC;
  SIGNAL and_dcpl_1127 : STD_LOGIC;
  SIGNAL and_dcpl_1130 : STD_LOGIC;
  SIGNAL and_dcpl_1141 : STD_LOGIC;
  SIGNAL and_dcpl_1145 : STD_LOGIC;
  SIGNAL and_dcpl_1151 : STD_LOGIC;
  SIGNAL and_dcpl_1152 : STD_LOGIC;
  SIGNAL or_tmp_1664 : STD_LOGIC;
  SIGNAL mux_tmp_2116 : STD_LOGIC;
  SIGNAL nand_tmp_99 : STD_LOGIC;
  SIGNAL mux_tmp_2119 : STD_LOGIC;
  SIGNAL or_tmp_1671 : STD_LOGIC;
  SIGNAL mux_tmp_2121 : STD_LOGIC;
  SIGNAL and_dcpl_1154 : STD_LOGIC;
  SIGNAL and_dcpl_1162 : STD_LOGIC;
  SIGNAL or_tmp_1690 : STD_LOGIC;
  SIGNAL mux_tmp_2153 : STD_LOGIC;
  SIGNAL or_dcpl_1178 : STD_LOGIC;
  SIGNAL mux_tmp_2176 : STD_LOGIC;
  SIGNAL or_dcpl_1180 : STD_LOGIC;
  SIGNAL or_dcpl_1181 : STD_LOGIC;
  SIGNAL or_dcpl_1183 : STD_LOGIC;
  SIGNAL or_dcpl_1184 : STD_LOGIC;
  SIGNAL or_dcpl_1186 : STD_LOGIC;
  SIGNAL or_dcpl_1187 : STD_LOGIC;
  SIGNAL or_dcpl_1188 : STD_LOGIC;
  SIGNAL or_dcpl_1189 : STD_LOGIC;
  SIGNAL and_dcpl_1193 : STD_LOGIC;
  SIGNAL and_dcpl_1194 : STD_LOGIC;
  SIGNAL and_dcpl_1195 : STD_LOGIC;
  SIGNAL or_dcpl_1195 : STD_LOGIC;
  SIGNAL or_dcpl_1196 : STD_LOGIC;
  SIGNAL or_dcpl_1198 : STD_LOGIC;
  SIGNAL or_dcpl_1199 : STD_LOGIC;
  SIGNAL or_dcpl_1201 : STD_LOGIC;
  SIGNAL or_dcpl_1203 : STD_LOGIC;
  SIGNAL or_dcpl_1209 : STD_LOGIC;
  SIGNAL and_dcpl_1199 : STD_LOGIC;
  SIGNAL nand_tmp_104 : STD_LOGIC;
  SIGNAL mux_tmp_2252 : STD_LOGIC;
  SIGNAL and_dcpl_1225 : STD_LOGIC;
  SIGNAL and_dcpl_1227 : STD_LOGIC;
  SIGNAL and_dcpl_1232 : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_nand_seb : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse
      : STD_LOGIC;
  SIGNAL RESHAPE_2D_TO_3D_LOOP_2_2_and_cse : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_i_4_0_sva_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_2_2_and_30_m1c : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_2_2_and_30_m1c_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_2_mx0 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1
      : STD_LOGIC_VECTOR (35 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_1_sva_1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_2_sva_1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_3_sva_1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_stg_2_0_sva_1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_stg_2_1_sva_1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_stg_2_2_sva_1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_stg_2_3_sva_1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_stg_1_0_sva_1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_stg_1_1_sva_1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_stg_1_2_sva_1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_stg_1_3_sva_1 : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_and_30_m1c : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_and_30_m1c_1 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_sva : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL input_0_0_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva : STD_LOGIC;
  SIGNAL TRANSPOSE_LAST_TWO_DIMS_LOOP_3_k_2_0_sva_1 : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_conc_1_1_1_0_svs_1
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_2_2_unequal_tmp_mx0w0 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_l_and_ssc : STD_LOGIC;
  SIGNAL reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd : STD_LOGIC;
  SIGNAL reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 : STD_LOGIC;
  SIGNAL and_336_ssc : STD_LOGIC;
  SIGNAL mux_856_ssc : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_59_39
      : STD_LOGIC_VECTOR (20 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_38_0
      : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL mux_851_ssc : STD_LOGIC;
  SIGNAL and_321_ssc : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_39 : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_38_35 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL mux_2100_ssc : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0 : STD_LOGIC;
  SIGNAL attention_abs_qelse_and_ssc : STD_LOGIC;
  SIGNAL attention_abs_4_qelse_and_ssc : STD_LOGIC;
  SIGNAL for_1_for_and_cse : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_and_cse : STD_LOGIC;
  SIGNAL input_and_cse : STD_LOGIC;
  SIGNAL and_1555_cse : STD_LOGIC;
  SIGNAL or_1769_cse : STD_LOGIC;
  SIGNAL or_1732_cse : STD_LOGIC;
  SIGNAL or_1770_cse : STD_LOGIC;
  SIGNAL reg_strm_out_rsci_iswt0_cse : STD_LOGIC;
  SIGNAL reg_strm_in_rsci_iswt0_cse : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_and_3_cse : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_and_6_cse : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_and_7_cse : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_and_8_cse : STD_LOGIC;
  SIGNAL and_1474_cse : STD_LOGIC;
  SIGNAL and_1559_cse : STD_LOGIC;
  SIGNAL mux_806_cse : STD_LOGIC;
  SIGNAL or_2249_cse : STD_LOGIC;
  SIGNAL and_1773_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_cse : STD_LOGIC;
  SIGNAL or_2456_cse : STD_LOGIC;
  SIGNAL and_1651_cse : STD_LOGIC;
  SIGNAL or_1907_cse : STD_LOGIC;
  SIGNAL nand_365_cse : STD_LOGIC;
  SIGNAL or_2480_cse : STD_LOGIC;
  SIGNAL or_2486_cse : STD_LOGIC;
  SIGNAL or_2742_cse : STD_LOGIC;
  SIGNAL or_2736_cse : STD_LOGIC;
  SIGNAL or_1880_cse : STD_LOGIC;
  SIGNAL mux_792_cse : STD_LOGIC;
  SIGNAL or_1983_cse : STD_LOGIC;
  SIGNAL or_2457_cse : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_and_28_cse : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_and_cse : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_44_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_mux_14_cse : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_mux_13_cse : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_mux_11_cse : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_mux_9_cse : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_mux_7_cse : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL nor_1239_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_weights_and_cse : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_36_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_weights_and_12_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_weights_and_24_cse : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_46_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_8_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_16_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_24_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_32_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_40_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_48_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_56_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_64_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_72_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_80_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_88_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_96_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_104_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_and_112_cse : STD_LOGIC;
  SIGNAL and_1455_cse : STD_LOGIC;
  SIGNAL nor_176_cse : STD_LOGIC;
  SIGNAL or_76_cse : STD_LOGIC;
  SIGNAL or_130_cse : STD_LOGIC;
  SIGNAL and_28_cse : STD_LOGIC;
  SIGNAL nor_1229_cse : STD_LOGIC;
  SIGNAL and_1771_cse : STD_LOGIC;
  SIGNAL and_1762_cse : STD_LOGIC;
  SIGNAL or_3185_cse : STD_LOGIC;
  SIGNAL nor_366_cse : STD_LOGIC;
  SIGNAL nand_197_cse : STD_LOGIC;
  SIGNAL or_2699_cse : STD_LOGIC;
  SIGNAL or_1848_cse : STD_LOGIC;
  SIGNAL or_133_cse : STD_LOGIC;
  SIGNAL nor_777_cse : STD_LOGIC;
  SIGNAL nor_973_cse : STD_LOGIC;
  SIGNAL and_37_cse : STD_LOGIC;
  SIGNAL or_361_cse : STD_LOGIC;
  SIGNAL or_362_cse : STD_LOGIC;
  SIGNAL and_1638_cse : STD_LOGIC;
  SIGNAL or_1985_cse : STD_LOGIC;
  SIGNAL or_1984_cse : STD_LOGIC;
  SIGNAL nor_749_cse : STD_LOGIC;
  SIGNAL or_2455_cse : STD_LOGIC;
  SIGNAL or_1197_cse : STD_LOGIC;
  SIGNAL or_822_cse : STD_LOGIC;
  SIGNAL or_2460_cse : STD_LOGIC;
  SIGNAL or_1879_cse : STD_LOGIC;
  SIGNAL nor_1026_cse : STD_LOGIC;
  SIGNAL or_270_cse : STD_LOGIC;
  SIGNAL or_1767_cse : STD_LOGIC;
  SIGNAL or_1772_cse : STD_LOGIC;
  SIGNAL nor_717_cse : STD_LOGIC;
  SIGNAL and_1572_cse : STD_LOGIC;
  SIGNAL or_1908_cse : STD_LOGIC;
  SIGNAL or_255_cse : STD_LOGIC;
  SIGNAL or_1851_cse : STD_LOGIC;
  SIGNAL or_1835_cse : STD_LOGIC;
  SIGNAL or_1867_cse : STD_LOGIC;
  SIGNAL or_1420_cse : STD_LOGIC;
  SIGNAL mux_623_cse : STD_LOGIC;
  SIGNAL mux_528_cse : STD_LOGIC;
  SIGNAL and_1570_cse : STD_LOGIC;
  SIGNAL or_750_cse : STD_LOGIC;
  SIGNAL or_619_cse : STD_LOGIC;
  SIGNAL or_790_cse : STD_LOGIC;
  SIGNAL nand_143_cse : STD_LOGIC;
  SIGNAL or_262_cse : STD_LOGIC;
  SIGNAL or_1435_cse : STD_LOGIC;
  SIGNAL or_806_cse : STD_LOGIC;
  SIGNAL or_1431_cse : STD_LOGIC;
  SIGNAL or_753_cse : STD_LOGIC;
  SIGNAL nor_992_cse : STD_LOGIC;
  SIGNAL or_2792_cse : STD_LOGIC;
  SIGNAL or_1795_cse : STD_LOGIC;
  SIGNAL nand_253_cse : STD_LOGIC;
  SIGNAL or_349_cse : STD_LOGIC;
  SIGNAL or_241_cse : STD_LOGIC;
  SIGNAL or_2451_cse : STD_LOGIC;
  SIGNAL nor_646_cse : STD_LOGIC;
  SIGNAL nand_129_cse : STD_LOGIC;
  SIGNAL or_3167_cse : STD_LOGIC;
  SIGNAL nor_354_cse : STD_LOGIC;
  SIGNAL nor_355_cse : STD_LOGIC;
  SIGNAL or_2395_cse : STD_LOGIC;
  SIGNAL nand_163_cse : STD_LOGIC;
  SIGNAL nand_240_cse : STD_LOGIC;
  SIGNAL nor_964_cse : STD_LOGIC;
  SIGNAL nand_263_cse : STD_LOGIC;
  SIGNAL or_2834_cse : STD_LOGIC;
  SIGNAL or_2797_cse : STD_LOGIC;
  SIGNAL nand_381_cse : STD_LOGIC;
  SIGNAL or_2029_cse : STD_LOGIC;
  SIGNAL nor_1106_cse : STD_LOGIC;
  SIGNAL nor_593_cse : STD_LOGIC;
  SIGNAL or_2500_cse : STD_LOGIC;
  SIGNAL or_2154_cse : STD_LOGIC;
  SIGNAL or_2739_cse : STD_LOGIC;
  SIGNAL or_3039_cse : STD_LOGIC;
  SIGNAL and_1782_cse : STD_LOGIC;
  SIGNAL or_3163_cse : STD_LOGIC;
  SIGNAL nor_305_cse : STD_LOGIC;
  SIGNAL or_2671_cse : STD_LOGIC;
  SIGNAL and_1790_cse : STD_LOGIC;
  SIGNAL mux_816_ssc : STD_LOGIC;
  SIGNAL reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd : STD_LOGIC;
  SIGNAL reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd_1 : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_i_and_ssc : STD_LOGIC;
  SIGNAL reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 : STD_LOGIC;
  SIGNAL reg_rms_norm_16_div_cmp_a_ftd : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL and_937_ssc : STD_LOGIC;
  SIGNAL nor_1324_seb : STD_LOGIC;
  SIGNAL CACHE_UPDATE_LOOP_3_k_and_ssc : STD_LOGIC;
  SIGNAL reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_17_16
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1 : STD_LOGIC;
  SIGNAL reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 : STD_LOGIC;
  SIGNAL for_for_and_13_ssc : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_or_cse : STD_LOGIC;
  SIGNAL mux_1639_cse : STD_LOGIC;
  SIGNAL mux_1551_cse : STD_LOGIC;
  SIGNAL or_2481_cse : STD_LOGIC;
  SIGNAL mux_1812_cse : STD_LOGIC;
  SIGNAL mux_1809_cse : STD_LOGIC;
  SIGNAL mux_2025_cse : STD_LOGIC;
  SIGNAL mux_2157_cse : STD_LOGIC;
  SIGNAL mux_958_cse : STD_LOGIC;
  SIGNAL and_1637_cse : STD_LOGIC;
  SIGNAL mux_2024_cse : STD_LOGIC;
  SIGNAL or_2717_cse : STD_LOGIC;
  SIGNAL mux_502_cse : STD_LOGIC;
  SIGNAL mux_304_cse : STD_LOGIC;
  SIGNAL mux_1522_cse : STD_LOGIC;
  SIGNAL or_3137_cse : STD_LOGIC;
  SIGNAL mux_624_cse : STD_LOGIC;
  SIGNAL nor_998_cse : STD_LOGIC;
  SIGNAL nand_50_cse : STD_LOGIC;
  SIGNAL mux_1074_cse : STD_LOGIC;
  SIGNAL mux_1089_cse : STD_LOGIC;
  SIGNAL mux_1087_cse : STD_LOGIC;
  SIGNAL mux_1084_cse : STD_LOGIC;
  SIGNAL mux_1309_cse : STD_LOGIC;
  SIGNAL mux_2092_cse : STD_LOGIC;
  SIGNAL and_1811_cse : STD_LOGIC;
  SIGNAL and_1781_cse : STD_LOGIC;
  SIGNAL mux_2139_cse : STD_LOGIC;
  SIGNAL or_2858_cse : STD_LOGIC;
  SIGNAL or_2856_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_and_4_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_weights_and_36_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_5_cse : STD_LOGIC;
  SIGNAL mux_1559_cse : STD_LOGIC;
  SIGNAL mux_1557_cse : STD_LOGIC;
  SIGNAL mux_1555_cse : STD_LOGIC;
  SIGNAL mux_1553_cse : STD_LOGIC;
  SIGNAL mux_1645_cse : STD_LOGIC;
  SIGNAL mux_1546_cse : STD_LOGIC;
  SIGNAL mux_2032_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_32_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_weights_and_48_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_63_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_65_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_67_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_69_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_71_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_73_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_75_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_77_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_79_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_81_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_83_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_85_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_87_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_89_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_91_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_93_cse : STD_LOGIC;
  SIGNAL output_and_16_cse : STD_LOGIC;
  SIGNAL mux_1122_cse : STD_LOGIC;
  SIGNAL mux_1125_cse : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c4 : STD_LOGIC;
  SIGNAL and_1191_rgt : STD_LOGIC;
  SIGNAL and_622_rgt : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_and_ssc : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_15
      : STD_LOGIC;
  SIGNAL mux_1132_cse : STD_LOGIC;
  SIGNAL CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_sdt : STD_LOGIC_VECTOR
      (19 DOWNTO 0);
  SIGNAL and_362_ssc : STD_LOGIC;
  SIGNAL TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_16_psp_1 : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL GEMM_3D_FLOAT_LOOP_4_acc_sdt_1 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_4_acc_13_sdt_1 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_acc_12_sdt_1 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL CACHE_UPDATE_LOOP_3_acc_sdt_1 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_sdt_1 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_0_0_0_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_2_0_3_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_3_0_0_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_3_0_1_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_3_0_2_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_dcpl_1233 : STD_LOGIC;
  SIGNAL attention_abs_qr_35_0_lpi_1_dfm_mx0w0 : STD_LOGIC_VECTOR (35 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva_mx0w0 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva_mx0w0 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva_mx0w0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c10 : STD_LOGIC;
  SIGNAL input_0_4_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c10 : STD_LOGIC;
  SIGNAL input_0_11_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c10 : STD_LOGIC;
  SIGNAL input_0_3_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL for_for_strm_in_tmp_sva_31_26 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL for_for_strm_in_tmp_sva_25_2 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c12 : STD_LOGIC;
  SIGNAL or_3212_tmp : STD_LOGIC;
  SIGNAL or_3213_tmp : STD_LOGIC;
  SIGNAL or_3214_tmp : STD_LOGIC;
  SIGNAL nand_303_tmp : STD_LOGIC;
  SIGNAL nand_304_tmp : STD_LOGIC;
  SIGNAL nand_305_tmp : STD_LOGIC;
  SIGNAL and_343_itm : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_mux1h_5_itm : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL and_404_itm : STD_LOGIC;
  SIGNAL and_416_itm : STD_LOGIC;
  SIGNAL and_428_itm : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_itm
      : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_itm
      : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_itm : STD_LOGIC_VECTOR
      (14 DOWNTO 0);
  SIGNAL and_615_itm : STD_LOGIC;
  SIGNAL and_633_itm : STD_LOGIC;
  SIGNAL and_654_itm : STD_LOGIC;
  SIGNAL and_648_itm : STD_LOGIC;
  SIGNAL and_642_itm : STD_LOGIC;
  SIGNAL and_636_itm : STD_LOGIC;
  SIGNAL and_629_itm : STD_LOGIC;
  SIGNAL and_639_itm : STD_LOGIC;
  SIGNAL and_645_itm : STD_LOGIC;
  SIGNAL and_651_itm : STD_LOGIC;
  SIGNAL and_657_itm : STD_LOGIC;
  SIGNAL nor_1144_itm : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm : STD_LOGIC_VECTOR
      (12 DOWNTO 0);
  SIGNAL and_1060_itm : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm
      : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm
      : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL mux_2256_itm : STD_LOGIC;
  SIGNAL mux_1147_itm : STD_LOGIC;
  SIGNAL mux_1177_itm : STD_LOGIC;
  SIGNAL mux_1197_itm : STD_LOGIC;
  SIGNAL CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_itm : STD_LOGIC_VECTOR
      (18 DOWNTO 0);
  SIGNAL and_dcpl_1248 : STD_LOGIC;
  SIGNAL z_out : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL and_dcpl_1261 : STD_LOGIC;
  SIGNAL z_out_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL and_dcpl_1273 : STD_LOGIC;
  SIGNAL z_out_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL and_dcpl_1294 : STD_LOGIC;
  SIGNAL z_out_3 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL z_out_4 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL z_out_5 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL and_dcpl_1363 : STD_LOGIC;
  SIGNAL and_dcpl_1371 : STD_LOGIC;
  SIGNAL and_dcpl_1379 : STD_LOGIC;
  SIGNAL and_dcpl_1385 : STD_LOGIC;
  SIGNAL z_out_9 : STD_LOGIC_VECTOR (59 DOWNTO 0);
  SIGNAL and_dcpl_1391 : STD_LOGIC;
  SIGNAL and_dcpl_1392 : STD_LOGIC;
  SIGNAL and_dcpl_1393 : STD_LOGIC;
  SIGNAL and_dcpl_1396 : STD_LOGIC;
  SIGNAL and_dcpl_1398 : STD_LOGIC;
  SIGNAL and_dcpl_1401 : STD_LOGIC;
  SIGNAL and_dcpl_1403 : STD_LOGIC;
  SIGNAL and_dcpl_1406 : STD_LOGIC;
  SIGNAL and_dcpl_1407 : STD_LOGIC;
  SIGNAL and_dcpl_1410 : STD_LOGIC;
  SIGNAL and_dcpl_1415 : STD_LOGIC;
  SIGNAL and_dcpl_1420 : STD_LOGIC;
  SIGNAL and_dcpl_1425 : STD_LOGIC;
  SIGNAL and_dcpl_1427 : STD_LOGIC;
  SIGNAL and_dcpl_1429 : STD_LOGIC;
  SIGNAL and_dcpl_1431 : STD_LOGIC;
  SIGNAL and_dcpl_1436 : STD_LOGIC;
  SIGNAL z_out_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_dcpl_1447 : STD_LOGIC;
  SIGNAL z_out_11 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL z_out_12 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL input_0_7_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_8_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_6_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_9_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_5_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_10_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_12_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_1_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_14_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_7_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_8_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_6_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_9_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_5_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_10_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_4_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_11_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_3_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_12_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_1_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_14_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL input_0_15_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_2_0_3_lpi_3 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_3_0_0_lpi_3 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_3_0_1_lpi_3 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_3_0_2_lpi_3 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_3_0_3_lpi_3 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_2_0_1_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_1_0_1_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_2_0_3_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_3_0_0_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_0_0_2_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_3_0_1_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_3_0_2_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_0_0_0_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_3_0_3_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_3 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_4 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_5 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_4 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_4 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_5 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_4 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_4 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_5 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_4 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_4 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_5 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_4 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL softmax_1_4_3_sum_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_0_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_1_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_2_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_3_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_2_and_29_ssc : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_and_34_ssc : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_and_29_ssc : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_and_34_ssc : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_mul_mut : STD_LOGIC_VECTOR (59 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_3_mul_mut : STD_LOGIC_VECTOR (59 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut : STD_LOGIC_VECTOR (60 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_mux1h_itm : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_mul_itm : STD_LOGIC_VECTOR (59 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mul_itm : STD_LOGIC_VECTOR (55 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mul_1_itm : STD_LOGIC_VECTOR (55 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm : STD_LOGIC_VECTOR (55 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mul_3_itm : STD_LOGIC_VECTOR (55 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_mux1h_itm : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_38_0 : STD_LOGIC_VECTOR (38 DOWNTO
      0);
  SIGNAL QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_38_0 : STD_LOGIC_VECTOR (38 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_7_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_8_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_6_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_9_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_5_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_10_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_4_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_11_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_12_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_13_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_14_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_0_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_15_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_7_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_8_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_6_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_9_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_5_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_10_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_4_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_11_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_12_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_13_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_14_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_0_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_15_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_7_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_8_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_6_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_9_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_5_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_10_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_4_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_11_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_12_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_13_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_14_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_0_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_15_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_7_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_15_0 : STD_LOGIC_VECTOR (15
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0 : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL output_0_7_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_7_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_8_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_8_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_6_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_6_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_9_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_9_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_5_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_5_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_10_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_10_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_4_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_4_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_11_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_11_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_3_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_3_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_12_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_12_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_2_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_2_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_13_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_13_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_1_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_14_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_14_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_0_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_0_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_15_lpi_3_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_15_lpi_3_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_7_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_8_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_6_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_9_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_5_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_10_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_4_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_11_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_3_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_12_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_2_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_13_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_1_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_14_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_0_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_15_lpi_4_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_7_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_8_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_6_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_9_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_5_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_10_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_4_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_11_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_3_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_12_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_2_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_13_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_1_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_14_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_0_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_15_sva_1_39_16 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_7_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_8_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_6_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_9_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_5_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_10_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_4_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_11_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_3_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_12_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_2_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_13_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_14_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_0_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL output_0_15_sva_2_15_0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48 : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16 : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_39_16 : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2_mx1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2_mx1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2_mx1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2_mx1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2_mx1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2_mx1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2_mx1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2_mx1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2_mx1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2_mx1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1_mx0w1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2_mx0w1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2_mx0w1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2_mx0w1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2_mx0w1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w0 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w3 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2_mx0w1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16_mx0w1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0_mx0w1 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL drf_output_sdt_2_sva_15_0_mx0w0 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL drf_output_sdt_3_sva_15_0_mx0w3 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL SOFTMAX_LOOP_5_mux_12_psp_mx0w0 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_conc_1_mut_71_48_mx0w0 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_3_conc_1_mut_71_48_mx0w3 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2 : STD_LOGIC_VECTOR (60 DOWNTO
      0);
  SIGNAL rms_norm_16_div_cmp_a_mx0c0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c9 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx2 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_abs_1_qr_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL softmax_1_4_3_sum_sva_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c0 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c2 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c3 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c5 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c7 : STD_LOGIC;
  SIGNAL for_for_strm_in_tmp_sva_31_2_mx0c1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c0 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c2 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c4 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c7 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c9 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c10 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c9 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx2 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c9 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c8 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c10 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c0 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c2 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c3 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c6 : STD_LOGIC;
  SIGNAL attention_abs_qr_35_0_lpi_1_dfm_mx0c1 : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_dfm_1_38_0_1 : STD_LOGIC_VECTOR
      (38 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c1 : STD_LOGIC;
  SIGNAL TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3 : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL CACHE_UPDATE_LOOP_3_k_2_0_sva_1_mx0c1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c2 : STD_LOGIC;
  SIGNAL attention_abs_2_mux_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_2_and_29_ssc_1 : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_and_34_ssc_1 : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_and_32_ssc_mx0w3 : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_nor_1_ssc_1 : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_and_33_ssc_1 : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_dfm_1_38_0_mx0w1 : STD_LOGIC_VECTOR
      (38 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16_mx0c1 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c0 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c2 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c3 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c8 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0_mx0w6 : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16_mx0c1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16_mx0c1 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48_mx0w2 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16_mx0w5 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_2 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1
      : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1
      : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1 :
      STD_LOGIC;
  SIGNAL RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1
      : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_4_sva_mx0w2 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_0_sva_mx0w3 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_5_sva_mx0w2 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_1_sva_mx0w3 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_6_sva_mx0w1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva_mx0w3 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_7_sva_mx0w1 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva_mx0w3 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1
      : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1
      : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1
      : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1
      : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c9 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx2 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx0c7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx0c7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c9 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx2 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx0c7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx0c7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx0c7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c9 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx2 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx0c7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_15_sdt_1 : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_sva_mx0w0 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva_mx0w0 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva_mx0w0 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva_mx0w0 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva_mx0w0 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva_mx0w0 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva_mx0w0 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva_mx0w0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1 : STD_LOGIC_VECTOR (38 DOWNTO
      0);
  SIGNAL SF_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_psp_sva_1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL CM_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_ctmp_sva_1 :
      STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8_mx1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL SOFTMAX_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_cse_sva_1
      : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL SOFTMAX_LOOP_4_acc_3_cse_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva_mx0w0 : STD_LOGIC;
  SIGNAL attention_abs_4_qr_35_0_lpi_1_dfm_mx0c1 : STD_LOGIC;
  SIGNAL attention_abs_5_qr_sva_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL attention_abs_6_mux_2 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_2_2_and_29_ssc_1 : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_and_34_ssc_1 : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_nor_1_ssc_1 : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_and_33_ssc_1 : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_nand_seb_1 : STD_LOGIC;
  SIGNAL output_0_15_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_0_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_14_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_1_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_13_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_2_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_12_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_3_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_11_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_4_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_10_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_5_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_9_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_6_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_8_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL output_0_7_lpi_4_39_16_mx1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_7_1 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_0_1 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_6_1 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_1_1 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_5_1 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_2_1 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_4_1 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_3_1 : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1 : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL attention_abs_3_qr_sva_38_0 : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL attention_abs_5_qr_sva_38_0 : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL attention_abs_7_qr_sva_38_0 : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL output_0_7_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_8_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_6_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_9_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_5_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_10_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_4_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_11_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_3_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_12_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_2_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_13_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_1_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_14_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_0_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL output_0_15_sva_2_29_16 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_39 :
      STD_LOGIC;
  SIGNAL attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_38_0
      : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL attention_abs_qr_35_0_lpi_1_dfm_35 : STD_LOGIC;
  SIGNAL attention_abs_qr_35_0_lpi_1_dfm_34_0 : STD_LOGIC_VECTOR (34 DOWNTO 0);
  SIGNAL attention_abs_4_qr_35_0_lpi_1_dfm_35 : STD_LOGIC;
  SIGNAL attention_abs_4_qr_35_0_lpi_1_dfm_34_0 : STD_LOGIC_VECTOR (34 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_conc_1_itm_11_0 : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_conc_3_itm_8_0 : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_or_3_ssc : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_or_1_ssc : STD_LOGIC;
  SIGNAL reg_rms_norm_16_div_cmp_b_ftd_1 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1 : STD_LOGIC_VECTOR
      (38 DOWNTO 0);
  SIGNAL reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd
      : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1
      : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2
      : STD_LOGIC;
  SIGNAL reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3
      : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_and_4_ssc : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_1 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_2 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_3 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_4 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_5 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_6 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_7 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd : STD_LOGIC_VECTOR (7
      DOWNTO 0);
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd : STD_LOGIC_VECTOR (7
      DOWNTO 0);
  SIGNAL and_581_ssc : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_nand_seb : STD_LOGIC;
  SIGNAL and_585_seb : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_1_ssc : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_or_1_cse : STD_LOGIC;
  SIGNAL rms_norm_16_variance_or_1_cse : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_and_14_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_and_13_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_and_16_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_and_15_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_and_18_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_and_17_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_and_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_and_1_cse : STD_LOGIC;
  SIGNAL nor_1053_cse : STD_LOGIC;
  SIGNAL nor_1044_cse : STD_LOGIC;
  SIGNAL nor_1045_cse : STD_LOGIC;
  SIGNAL nor_1138_m1c : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_47_40
      : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL reg_rms_norm_16_div_cmp_a_ftd_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_8_seb : STD_LOGIC;
  SIGNAL or_1667_ssc : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_39 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_38_0 : STD_LOGIC_VECTOR
      (38 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_7 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_6 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_5 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_4 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_3 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_2 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_1 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_0 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_7 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_6 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_5 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_4 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_3 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_2 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_1 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_0 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_7 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_6 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_5 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_4 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_3 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_2 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_1 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_39 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_38_0 : STD_LOGIC_VECTOR
      (38 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0 : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_or_2_ssc : STD_LOGIC;
  SIGNAL nor_1314_cse : STD_LOGIC;
  SIGNAL mux_1513_cse : STD_LOGIC;
  SIGNAL CACHE_UPDATE_LOOP_3_or_cse : STD_LOGIC;
  SIGNAL CACHE_UPDATE_LOOP_3_or_1_cse : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_or_5_cse : STD_LOGIC;
  SIGNAL compute_sqrt_for_i_and_2_cse : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_and_31_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1 : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_hidden_states_and_3_ssc : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_hidden_states_0_7_sva_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_hidden_states_and_2_ssc : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_hidden_states_0_8_sva_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_hidden_states_and_1_ssc : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_hidden_states_0_6_sva_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_hidden_states_and_ssc : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_quantized_hidden_states_0_9_sva_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_15 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_14_12 : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_11_9 : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_8 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 :
      STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 :
      STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL nor_1228_ssc : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_and_5_ssc : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_0 : STD_LOGIC;
  SIGNAL input_0_13_sva_1_39 : STD_LOGIC;
  SIGNAL input_0_13_sva_1_38_0 : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_and_29_ssc : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_cse : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_cse : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse : STD_LOGIC;
  SIGNAL and_474_rgt : STD_LOGIC;
  SIGNAL and_476_rgt : STD_LOGIC;
  SIGNAL and_480_rgt : STD_LOGIC;
  SIGNAL for_for_and_14_rgt : STD_LOGIC;
  SIGNAL for_for_and_15_rgt : STD_LOGIC;
  SIGNAL for_for_and_16_rgt : STD_LOGIC;
  SIGNAL for_for_and_17_rgt : STD_LOGIC;
  SIGNAL and_485_rgt : STD_LOGIC;
  SIGNAL and_486_rgt : STD_LOGIC;
  SIGNAL for_for_or_1_rgt : STD_LOGIC;
  SIGNAL and_745_ssc : STD_LOGIC;
  SIGNAL input_0_13_sva_2_39 : STD_LOGIC;
  SIGNAL input_0_13_sva_2_38_0 : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 :
      STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL attention_abs_qr_35_0_lpi_1_dfm_mx1_35 : STD_LOGIC;
  SIGNAL attention_abs_qr_35_0_lpi_1_dfm_mx1_34_1 : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_0 : STD_LOGIC;
  SIGNAL and_303_ssc : STD_LOGIC;
  SIGNAL compute_sqrt_guess_or_1_ssc : STD_LOGIC;
  SIGNAL and_315_ssc : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_34 : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_33_0 : STD_LOGIC_VECTOR (33
      DOWNTO 0);
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_and_ssc : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39 : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0 : STD_LOGIC_VECTOR
      (38 DOWNTO 0);
  SIGNAL compute_sqrt_guess_and_ssc : STD_LOGIC;
  SIGNAL compute_sqrt_guess_sva_34 : STD_LOGIC;
  SIGNAL compute_sqrt_guess_sva_33_0 : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL compute_sqrt_1_guess_and_ssc : STD_LOGIC;
  SIGNAL compute_sqrt_1_guess_sva_34 : STD_LOGIC;
  SIGNAL compute_sqrt_1_guess_sva_33_0 : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_or_11_cse : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_or_12_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_25_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_27_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_29_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_or_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_or_17_cse : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_i_and_9_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_and_91_cse : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_l_or_2_cse : STD_LOGIC;
  SIGNAL input_0_2_sva_1_39 : STD_LOGIC;
  SIGNAL input_0_2_sva_1_38_0 : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8
      : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL and_699_ssc : STD_LOGIC;
  SIGNAL input_0_2_sva_2_39 : STD_LOGIC;
  SIGNAL input_0_2_sva_2_38_0 : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 :
      STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_and_2_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_26_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_28_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_30_cse : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_and_4_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_re_and_29_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_and_65_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_and_95_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_and_30_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_weights_and_52_cse : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_ftd : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL and_1055_ssc : STD_LOGIC;
  SIGNAL and_1059_ssc : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_and_30_ssc : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL output_0_1_lpi_3_15_8 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL output_0_1_sva_2_15_8 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_proj_and_23_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_ftd : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL strm_out_rsci_idat_17_10 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL operator_80_48_true_AC_TRN_AC_WRAP_operator_80_48_true_AC_TRN_AC_WRAP_slc_SOFTMAX_LOOP_4_sqr_56_1_itm_slc
      : STD_LOGIC;
  SIGNAL reg_QUANTIZE_ACTIVATION_LOOP_3_quantized_value_slc_63_32_cse_slc : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL reg_RMS_NORM_LOOP_1_1_slc_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_mul_55_16_cse_1_slc
      : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL nand_302_cse : STD_LOGIC;
  SIGNAL RESHAPE_2D_TO_3D_LOOP_3_1_mux_13_cse : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_23_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_24_cse : STD_LOGIC;
  SIGNAL ATTN_2D_LOOP_3_mux_16_itm : STD_LOGIC;
  SIGNAL ATTN_2D_LOOP_3_mux_17_itm : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_nand_itm : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_5_itm : STD_LOGIC;
  SIGNAL mux_1512_itm : STD_LOGIC;
  SIGNAL and_1034_itm : STD_LOGIC;
  SIGNAL mux_1966_itm : STD_LOGIC;
  SIGNAL and_1037_itm : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm
      : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm
      : STD_LOGIC;
  SIGNAL mux_1079_itm : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_or_4_itm : STD_LOGIC;
  SIGNAL compute_sqrt_1_for_acc_1_itm_40_1_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL compute_sqrt_for_acc_1_itm_40_1_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL QUANTIZE_ACTIVATION_LOOP_2_acc_4_itm_40_1 : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_itm_40_1 : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1 : STD_LOGIC;
  SIGNAL CACHE_UPDATE_LOOP_2_1_acc_2_itm_2_1 : STD_LOGIC;
  SIGNAL attention_max_attn_fixed_t_1_acc_1_itm_40_1 : STD_LOGIC;
  SIGNAL CACHE_UPDATE_LOOP_2_acc_2_itm_2_1 : STD_LOGIC;
  SIGNAL SOFTMAX_LOOP_3_acc_3_itm_40_1 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_1 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_2 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_3 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_4 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_5 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_6 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_7 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_8 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_1 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_2 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_3 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_4 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_5 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_6 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_7 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_8 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_1 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_2 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_3 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_4 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_5 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_6 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_7 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_8 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_and_ssc : STD_LOGIC;
  SIGNAL reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd : STD_LOGIC;
  SIGNAL reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1 : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_ssc : STD_LOGIC;
  SIGNAL reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd : STD_LOGIC;
  SIGNAL reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 : STD_LOGIC;
  SIGNAL reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_and_ssc : STD_LOGIC;
  SIGNAL reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd : STD_LOGIC;
  SIGNAL reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_1_i_and_ssc : STD_LOGIC;
  SIGNAL reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd : STD_LOGIC;
  SIGNAL reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_1_i_and_ssc : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_k_and_ssc : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_and_18_ssc : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1 : STD_LOGIC_VECTOR
      (12 DOWNTO 0);
  SIGNAL reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd : STD_LOGIC;
  SIGNAL reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1 : STD_LOGIC;
  SIGNAL reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2 : STD_LOGIC;
  SIGNAL reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3 : STD_LOGIC;
  SIGNAL reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4 : STD_LOGIC;
  SIGNAL reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5 : STD_LOGIC;
  SIGNAL reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6 : STD_LOGIC;
  SIGNAL reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_and_17_ssc : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_0 : STD_LOGIC;
  SIGNAL and_1042_ssc : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_and_16_ssc : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 :
      STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_nor_seb : STD_LOGIC;
  SIGNAL and_1062_ssc : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_and_19_ssc : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_0 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_and_37_cse : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_and_25_cse : STD_LOGIC;
  SIGNAL input_and_28_cse : STD_LOGIC;
  SIGNAL output_and_64_cse : STD_LOGIC;
  SIGNAL and_339_ssc : STD_LOGIC;
  SIGNAL SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_39 : STD_LOGIC;
  SIGNAL SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_38_0 : STD_LOGIC_VECTOR (38 DOWNTO
      0);
  SIGNAL and_329_ssc : STD_LOGIC;
  SIGNAL and_334_ssc : STD_LOGIC;
  SIGNAL SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_55 : STD_LOGIC;
  SIGNAL SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_54_16 : STD_LOGIC_VECTOR (38 DOWNTO
      0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_1
      : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_0
      : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_15_13 : STD_LOGIC_VECTOR (2
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0 : STD_LOGIC_VECTOR (12
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_15_8 : STD_LOGIC_VECTOR (7
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_15_8 : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_15_13 : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0 : STD_LOGIC_VECTOR
      (12 DOWNTO 0);
  SIGNAL reg_rms_norm_16_div_cmp_b_ftd_59_38 : STD_LOGIC_VECTOR (21 DOWNTO 0);
  SIGNAL reg_rms_norm_16_div_cmp_b_ftd_37_0 : STD_LOGIC_VECTOR (37 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_39
      : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_38
      : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_37
      : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_36
      : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_35
      : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_34
      : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_33
      : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_32
      : STD_LOGIC;
  SIGNAL reg_rms_norm_16_div_cmp_a_ftd_1_7 : STD_LOGIC;
  SIGNAL reg_rms_norm_16_div_cmp_a_ftd_1_6 : STD_LOGIC;
  SIGNAL reg_rms_norm_16_div_cmp_a_ftd_1_5 : STD_LOGIC;
  SIGNAL reg_rms_norm_16_div_cmp_a_ftd_1_4 : STD_LOGIC;
  SIGNAL reg_rms_norm_16_div_cmp_a_ftd_1_3 : STD_LOGIC;
  SIGNAL reg_rms_norm_16_div_cmp_a_ftd_1_2 : STD_LOGIC;
  SIGNAL reg_rms_norm_16_div_cmp_a_ftd_1_1 : STD_LOGIC;
  SIGNAL reg_rms_norm_16_div_cmp_a_ftd_1_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_7 : STD_LOGIC;
  SIGNAL RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_6 : STD_LOGIC;
  SIGNAL RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_5 : STD_LOGIC;
  SIGNAL RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_4 : STD_LOGIC;
  SIGNAL RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_3 : STD_LOGIC;
  SIGNAL RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_2 : STD_LOGIC;
  SIGNAL RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_1 : STD_LOGIC;
  SIGNAL RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_13
      : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_12_8 :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_8 : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_13 : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0 : STD_LOGIC_VECTOR (12 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_13 : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_12_8 : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_1_or_ssc : STD_LOGIC;
  SIGNAL and_1908_cse : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1 : STD_LOGIC;
  SIGNAL reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0
      : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_1
      : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_0
      : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_0 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd :
      STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_1
      : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_2
      : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_3
      : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_4
      : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_5
      : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_6
      : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_7
      : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd :
      STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_1
      : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_2
      : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_3
      : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_4
      : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_5
      : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_6
      : STD_LOGIC;
  SIGNAL reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_7
      : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_1 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_2 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_3 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_4 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_5 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_6 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_7 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1 : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_0 : STD_LOGIC;
  SIGNAL output_0_1_lpi_3_7 : STD_LOGIC;
  SIGNAL output_0_1_lpi_3_6 : STD_LOGIC;
  SIGNAL output_0_1_lpi_3_5 : STD_LOGIC;
  SIGNAL output_0_1_lpi_3_4 : STD_LOGIC;
  SIGNAL output_0_1_lpi_3_3 : STD_LOGIC;
  SIGNAL output_0_1_lpi_3_2 : STD_LOGIC;
  SIGNAL output_0_1_lpi_3_1 : STD_LOGIC;
  SIGNAL output_0_1_lpi_3_0 : STD_LOGIC;
  SIGNAL output_0_1_sva_2_7 : STD_LOGIC;
  SIGNAL output_0_1_sva_2_6 : STD_LOGIC;
  SIGNAL output_0_1_sva_2_5 : STD_LOGIC;
  SIGNAL output_0_1_sva_2_4 : STD_LOGIC;
  SIGNAL output_0_1_sva_2_3 : STD_LOGIC;
  SIGNAL output_0_1_sva_2_2 : STD_LOGIC;
  SIGNAL output_0_1_sva_2_1 : STD_LOGIC;
  SIGNAL output_0_1_sva_2_0 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_7 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_6 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_5 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_4 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_3 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_2 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_1 : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_0 : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_7_cse : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_8_cse : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_9_cse : STD_LOGIC;
  SIGNAL compute_sqrt_for_i_and_cse : STD_LOGIC;
  SIGNAL compute_sqrt_for_i_and_4_cse : STD_LOGIC;
  SIGNAL compute_sqrt_for_i_and_5_cse : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_1 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_2 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_3 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_4 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_5 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_6 : STD_LOGIC;
  SIGNAL reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_7 : STD_LOGIC;
  SIGNAL strm_out_rsci_idat_9 : STD_LOGIC;
  SIGNAL strm_out_rsci_idat_8 : STD_LOGIC;
  SIGNAL strm_out_rsci_idat_7 : STD_LOGIC;
  SIGNAL strm_out_rsci_idat_6 : STD_LOGIC;
  SIGNAL strm_out_rsci_idat_5 : STD_LOGIC;
  SIGNAL strm_out_rsci_idat_4 : STD_LOGIC;
  SIGNAL strm_out_rsci_idat_3 : STD_LOGIC;
  SIGNAL strm_out_rsci_idat_2 : STD_LOGIC;
  SIGNAL z_out_13_71_28 : STD_LOGIC_VECTOR (43 DOWNTO 0);
  SIGNAL acc_3_cse_40_1 : STD_LOGIC_VECTOR (39 DOWNTO 0);

  SIGNAL mux_778_nl : STD_LOGIC;
  SIGNAL mux_777_nl : STD_LOGIC;
  SIGNAL mux_776_nl : STD_LOGIC;
  SIGNAL mux_775_nl : STD_LOGIC;
  SIGNAL and_1481_nl : STD_LOGIC;
  SIGNAL mux_774_nl : STD_LOGIC;
  SIGNAL or_1677_nl : STD_LOGIC;
  SIGNAL mux_773_nl : STD_LOGIC;
  SIGNAL or_1676_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_31_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_32_nl : STD_LOGIC;
  SIGNAL mux_786_nl : STD_LOGIC;
  SIGNAL mux_785_nl : STD_LOGIC;
  SIGNAL mux_784_nl : STD_LOGIC;
  SIGNAL mux_783_nl : STD_LOGIC;
  SIGNAL mux_782_nl : STD_LOGIC;
  SIGNAL mux_781_nl : STD_LOGIC;
  SIGNAL nor_728_nl : STD_LOGIC;
  SIGNAL mux_780_nl : STD_LOGIC;
  SIGNAL mux_779_nl : STD_LOGIC;
  SIGNAL and_1383_nl : STD_LOGIC;
  SIGNAL and_1485_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_32_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_4_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_34_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_6_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_30_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_2_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_40_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_12_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_42_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_14_nl : STD_LOGIC;
  SIGNAL and_259_nl : STD_LOGIC;
  SIGNAL mux_789_nl : STD_LOGIC;
  SIGNAL and_267_nl : STD_LOGIC;
  SIGNAL mux_797_nl : STD_LOGIC;
  SIGNAL mux_796_nl : STD_LOGIC;
  SIGNAL mux_795_nl : STD_LOGIC;
  SIGNAL mux_794_nl : STD_LOGIC;
  SIGNAL mux_793_nl : STD_LOGIC;
  SIGNAL or_1734_nl : STD_LOGIC;
  SIGNAL mux_791_nl : STD_LOGIC;
  SIGNAL nand_307_nl : STD_LOGIC;
  SIGNAL mux_790_nl : STD_LOGIC;
  SIGNAL nand_308_nl : STD_LOGIC;
  SIGNAL nand_309_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_38_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_10_nl : STD_LOGIC;
  SIGNAL mux_804_nl : STD_LOGIC;
  SIGNAL mux_803_nl : STD_LOGIC;
  SIGNAL mux_802_nl : STD_LOGIC;
  SIGNAL mux_801_nl : STD_LOGIC;
  SIGNAL and_274_nl : STD_LOGIC;
  SIGNAL mux_800_nl : STD_LOGIC;
  SIGNAL mux_799_nl : STD_LOGIC;
  SIGNAL nor_271_nl : STD_LOGIC;
  SIGNAL mux_815_nl : STD_LOGIC;
  SIGNAL mux_814_nl : STD_LOGIC;
  SIGNAL or_1775_nl : STD_LOGIC;
  SIGNAL or_1774_nl : STD_LOGIC;
  SIGNAL mux_813_nl : STD_LOGIC;
  SIGNAL mux_812_nl : STD_LOGIC;
  SIGNAL or_1771_nl : STD_LOGIC;
  SIGNAL mux_811_nl : STD_LOGIC;
  SIGNAL nand_41_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_nl : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL not_4947_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_1_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_2_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_3_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_4_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_5_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_6_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_7_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_8_nl : STD_LOGIC;
  SIGNAL mux_838_nl : STD_LOGIC;
  SIGNAL mux_850_nl : STD_LOGIC;
  SIGNAL mux_849_nl : STD_LOGIC;
  SIGNAL or_1803_nl : STD_LOGIC;
  SIGNAL mux_848_nl : STD_LOGIC;
  SIGNAL mux_847_nl : STD_LOGIC;
  SIGNAL mux_846_nl : STD_LOGIC;
  SIGNAL or_1802_nl : STD_LOGIC;
  SIGNAL mux_845_nl : STD_LOGIC;
  SIGNAL or_1799_nl : STD_LOGIC;
  SIGNAL mux_844_nl : STD_LOGIC;
  SIGNAL mux_843_nl : STD_LOGIC;
  SIGNAL mux_842_nl : STD_LOGIC;
  SIGNAL or_1798_nl : STD_LOGIC;
  SIGNAL mux_840_nl : STD_LOGIC;
  SIGNAL or_1792_nl : STD_LOGIC;
  SIGNAL mux_853_nl : STD_LOGIC;
  SIGNAL nor_977_nl : STD_LOGIC;
  SIGNAL and_1562_nl : STD_LOGIC;
  SIGNAL mux_852_nl : STD_LOGIC;
  SIGNAL and_1561_nl : STD_LOGIC;
  SIGNAL rms_norm_16_mux1h_nl : STD_LOGIC;
  SIGNAL rms_norm_16_mux1h_9_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_not_1_nl : STD_LOGIC;
  SIGNAL mux_854_nl : STD_LOGIC;
  SIGNAL SOFTMAX_LOOP_5_mux_24_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_mux1h_2_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_not_nl : STD_LOGIC;
  SIGNAL nor_979_nl : STD_LOGIC;
  SIGNAL mux_855_nl : STD_LOGIC;
  SIGNAL or_1812_nl : STD_LOGIC;
  SIGNAL and_1564_nl : STD_LOGIC;
  SIGNAL mux_861_nl : STD_LOGIC;
  SIGNAL mux_860_nl : STD_LOGIC;
  SIGNAL mux_859_nl : STD_LOGIC;
  SIGNAL mux_862_nl : STD_LOGIC;
  SIGNAL mux_864_nl : STD_LOGIC;
  SIGNAL mux_863_nl : STD_LOGIC;
  SIGNAL rms_norm_16_mux1h_10_nl : STD_LOGIC;
  SIGNAL rms_norm_16_mux1h_6_nl : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL rms_norm_16_not_nl : STD_LOGIC;
  SIGNAL rms_norm_16_mux1h_7_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL rms_norm_16_not_1_nl : STD_LOGIC;
  SIGNAL rms_norm_16_mux1h_11_nl : STD_LOGIC;
  SIGNAL rms_norm_16_mux1h_13_nl : STD_LOGIC;
  SIGNAL rms_norm_16_mux1h_14_nl : STD_LOGIC;
  SIGNAL rms_norm_16_mux1h_15_nl : STD_LOGIC;
  SIGNAL rms_norm_16_mux1h_16_nl : STD_LOGIC;
  SIGNAL rms_norm_16_mux1h_17_nl : STD_LOGIC;
  SIGNAL rms_norm_16_mux1h_18_nl : STD_LOGIC;
  SIGNAL rms_norm_16_mux1h_19_nl : STD_LOGIC;
  SIGNAL mux_874_nl : STD_LOGIC;
  SIGNAL mux_873_nl : STD_LOGIC;
  SIGNAL nor_907_nl : STD_LOGIC;
  SIGNAL mux_872_nl : STD_LOGIC;
  SIGNAL mux_871_nl : STD_LOGIC;
  SIGNAL mux_870_nl : STD_LOGIC;
  SIGNAL or_85_nl : STD_LOGIC;
  SIGNAL mux_878_nl : STD_LOGIC;
  SIGNAL mux_877_nl : STD_LOGIC;
  SIGNAL mux_876_nl : STD_LOGIC;
  SIGNAL nor_294_nl : STD_LOGIC;
  SIGNAL mux_882_nl : STD_LOGIC;
  SIGNAL mux_881_nl : STD_LOGIC;
  SIGNAL mux_880_nl : STD_LOGIC;
  SIGNAL or_1840_nl : STD_LOGIC;
  SIGNAL mux_886_nl : STD_LOGIC;
  SIGNAL mux_885_nl : STD_LOGIC;
  SIGNAL mux_884_nl : STD_LOGIC;
  SIGNAL nor_301_nl : STD_LOGIC;
  SIGNAL mux_902_nl : STD_LOGIC;
  SIGNAL mux_901_nl : STD_LOGIC;
  SIGNAL or_1857_nl : STD_LOGIC;
  SIGNAL mux_900_nl : STD_LOGIC;
  SIGNAL mux_899_nl : STD_LOGIC;
  SIGNAL mux_898_nl : STD_LOGIC;
  SIGNAL mux_897_nl : STD_LOGIC;
  SIGNAL nor_980_nl : STD_LOGIC;
  SIGNAL nor_981_nl : STD_LOGIC;
  SIGNAL or_1854_nl : STD_LOGIC;
  SIGNAL mux_896_nl : STD_LOGIC;
  SIGNAL or_1853_nl : STD_LOGIC;
  SIGNAL mux_895_nl : STD_LOGIC;
  SIGNAL mux_894_nl : STD_LOGIC;
  SIGNAL and_380_nl : STD_LOGIC;
  SIGNAL mux_893_nl : STD_LOGIC;
  SIGNAL mux_892_nl : STD_LOGIC;
  SIGNAL mux_891_nl : STD_LOGIC;
  SIGNAL nand_316_nl : STD_LOGIC;
  SIGNAL or_1849_nl : STD_LOGIC;
  SIGNAL mux_890_nl : STD_LOGIC;
  SIGNAL mux_889_nl : STD_LOGIC;
  SIGNAL mux_888_nl : STD_LOGIC;
  SIGNAL or_1847_nl : STD_LOGIC;
  SIGNAL mux_887_nl : STD_LOGIC;
  SIGNAL or_1846_nl : STD_LOGIC;
  SIGNAL or_1845_nl : STD_LOGIC;
  SIGNAL mux_905_nl : STD_LOGIC;
  SIGNAL or_3156_nl : STD_LOGIC;
  SIGNAL or_3157_nl : STD_LOGIC;
  SIGNAL mux_948_nl : STD_LOGIC;
  SIGNAL nor_985_nl : STD_LOGIC;
  SIGNAL mux_947_nl : STD_LOGIC;
  SIGNAL and_1566_nl : STD_LOGIC;
  SIGNAL nor_986_nl : STD_LOGIC;
  SIGNAL mux_946_nl : STD_LOGIC;
  SIGNAL mux_945_nl : STD_LOGIC;
  SIGNAL mux_944_nl : STD_LOGIC;
  SIGNAL mux_943_nl : STD_LOGIC;
  SIGNAL mux_942_nl : STD_LOGIC;
  SIGNAL mux_941_nl : STD_LOGIC;
  SIGNAL mux_940_nl : STD_LOGIC;
  SIGNAL mux_939_nl : STD_LOGIC;
  SIGNAL mux_938_nl : STD_LOGIC;
  SIGNAL mux_935_nl : STD_LOGIC;
  SIGNAL mux_934_nl : STD_LOGIC;
  SIGNAL mux_933_nl : STD_LOGIC;
  SIGNAL mux_932_nl : STD_LOGIC;
  SIGNAL mux_931_nl : STD_LOGIC;
  SIGNAL mux_930_nl : STD_LOGIC;
  SIGNAL mux_929_nl : STD_LOGIC;
  SIGNAL mux_928_nl : STD_LOGIC;
  SIGNAL mux_926_nl : STD_LOGIC;
  SIGNAL mux_925_nl : STD_LOGIC;
  SIGNAL mux_924_nl : STD_LOGIC;
  SIGNAL mux_923_nl : STD_LOGIC;
  SIGNAL mux_920_nl : STD_LOGIC;
  SIGNAL mux_918_nl : STD_LOGIC;
  SIGNAL mux_917_nl : STD_LOGIC;
  SIGNAL mux_914_nl : STD_LOGIC;
  SIGNAL mux_913_nl : STD_LOGIC;
  SIGNAL mux_912_nl : STD_LOGIC;
  SIGNAL mux_911_nl : STD_LOGIC;
  SIGNAL mux_907_nl : STD_LOGIC;
  SIGNAL rms_norm_16_variance_mux1h_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_mux_17_nl : STD_LOGIC;
  SIGNAL rms_norm_16_variance_mux1h_1_nl : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_mux_24_nl : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL mux_952_nl : STD_LOGIC;
  SIGNAL nor_990_nl : STD_LOGIC;
  SIGNAL mux_951_nl : STD_LOGIC;
  SIGNAL or_1890_nl : STD_LOGIC;
  SIGNAL or_1889_nl : STD_LOGIC;
  SIGNAL mux_950_nl : STD_LOGIC;
  SIGNAL or_3158_nl : STD_LOGIC;
  SIGNAL nand_318_nl : STD_LOGIC;
  SIGNAL and_1568_nl : STD_LOGIC;
  SIGNAL mux_949_nl : STD_LOGIC;
  SIGNAL nor_988_nl : STD_LOGIC;
  SIGNAL nor_989_nl : STD_LOGIC;
  SIGNAL mux_985_nl : STD_LOGIC;
  SIGNAL nand_47_nl : STD_LOGIC;
  SIGNAL mux_2236_nl : STD_LOGIC;
  SIGNAL or_3206_nl : STD_LOGIC;
  SIGNAL or_3207_nl : STD_LOGIC;
  SIGNAL mux_981_nl : STD_LOGIC;
  SIGNAL or_3159_nl : STD_LOGIC;
  SIGNAL mux_980_nl : STD_LOGIC;
  SIGNAL mux_979_nl : STD_LOGIC;
  SIGNAL mux_978_nl : STD_LOGIC;
  SIGNAL or_1923_nl : STD_LOGIC;
  SIGNAL or_1922_nl : STD_LOGIC;
  SIGNAL or_1920_nl : STD_LOGIC;
  SIGNAL mux_977_nl : STD_LOGIC;
  SIGNAL or_1919_nl : STD_LOGIC;
  SIGNAL or_1918_nl : STD_LOGIC;
  SIGNAL or_3160_nl : STD_LOGIC;
  SIGNAL mux_976_nl : STD_LOGIC;
  SIGNAL or_1916_nl : STD_LOGIC;
  SIGNAL nand_321_nl : STD_LOGIC;
  SIGNAL mux_974_nl : STD_LOGIC;
  SIGNAL mux_973_nl : STD_LOGIC;
  SIGNAL mux_972_nl : STD_LOGIC;
  SIGNAL mux_971_nl : STD_LOGIC;
  SIGNAL mux_970_nl : STD_LOGIC;
  SIGNAL mux_969_nl : STD_LOGIC;
  SIGNAL nor_991_nl : STD_LOGIC;
  SIGNAL mux_966_nl : STD_LOGIC;
  SIGNAL mux_965_nl : STD_LOGIC;
  SIGNAL mux_964_nl : STD_LOGIC;
  SIGNAL mux_963_nl : STD_LOGIC;
  SIGNAL mux_961_nl : STD_LOGIC;
  SIGNAL nand_319_nl : STD_LOGIC;
  SIGNAL mux_959_nl : STD_LOGIC;
  SIGNAL mux_957_nl : STD_LOGIC;
  SIGNAL or_1901_nl : STD_LOGIC;
  SIGNAL or_1899_nl : STD_LOGIC;
  SIGNAL nand_46_nl : STD_LOGIC;
  SIGNAL mux_956_nl : STD_LOGIC;
  SIGNAL mux_955_nl : STD_LOGIC;
  SIGNAL mux_954_nl : STD_LOGIC;
  SIGNAL or_1898_nl : STD_LOGIC;
  SIGNAL or_1895_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux_nl
      : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_8_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_9_nl : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_1_nl
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux_nl : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL and_1238_nl : STD_LOGIC;
  SIGNAL nor_1322_nl : STD_LOGIC;
  SIGNAL mux_2232_nl : STD_LOGIC;
  SIGNAL mux_2231_nl : STD_LOGIC;
  SIGNAL mux_2230_nl : STD_LOGIC;
  SIGNAL and_426_nl : STD_LOGIC;
  SIGNAL mux_984_nl : STD_LOGIC;
  SIGNAL mux_983_nl : STD_LOGIC;
  SIGNAL nor_996_nl : STD_LOGIC;
  SIGNAL mux_982_nl : STD_LOGIC;
  SIGNAL compute_sqrt_for_i_mux1h_nl : STD_LOGIC;
  SIGNAL mux_2229_nl : STD_LOGIC;
  SIGNAL mux_2228_nl : STD_LOGIC;
  SIGNAL mux_2227_nl : STD_LOGIC;
  SIGNAL nor_1311_nl : STD_LOGIC;
  SIGNAL compute_sqrt_for_i_nand_1_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL compute_sqrt_for_i_mux1h_1_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_not_2_nl : STD_LOGIC;
  SIGNAL compute_sqrt_for_i_mux1h_2_nl : STD_LOGIC;
  SIGNAL compute_sqrt_for_i_or_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_1_and_nl : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL INIT_2D_MEM_LOOP_2_1_mux1h_nl : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_37_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_69_nl : STD_LOGIC_VECTOR (22 DOWNTO 0);
  SIGNAL nor_1225_nl : STD_LOGIC;
  SIGNAL mux_2081_nl : STD_LOGIC;
  SIGNAL mux_2080_nl : STD_LOGIC;
  SIGNAL nand_373_nl : STD_LOGIC;
  SIGNAL mux_2079_nl : STD_LOGIC;
  SIGNAL nor_576_nl : STD_LOGIC;
  SIGNAL or_2777_nl : STD_LOGIC;
  SIGNAL mux_2077_nl : STD_LOGIC;
  SIGNAL or_2775_nl : STD_LOGIC;
  SIGNAL and_1110_nl : STD_LOGIC;
  SIGNAL and_1115_nl : STD_LOGIC;
  SIGNAL nor_1323_nl : STD_LOGIC;
  SIGNAL mux_2076_nl : STD_LOGIC;
  SIGNAL nand_96_nl : STD_LOGIC;
  SIGNAL mux_2075_nl : STD_LOGIC;
  SIGNAL mux_2074_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_mux_17_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL SOFTMAX_LOOP_4_x_acc_2_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL SOFTMAX_LOOP_4_x_mux_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_mux_18_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL mux_1063_nl : STD_LOGIC;
  SIGNAL mux_1062_nl : STD_LOGIC;
  SIGNAL mux_1061_nl : STD_LOGIC;
  SIGNAL mux_1060_nl : STD_LOGIC;
  SIGNAL mux_1059_nl : STD_LOGIC;
  SIGNAL mux_1058_nl : STD_LOGIC;
  SIGNAL mux_1057_nl : STD_LOGIC;
  SIGNAL mux_1056_nl : STD_LOGIC;
  SIGNAL mux_1055_nl : STD_LOGIC;
  SIGNAL mux_1054_nl : STD_LOGIC;
  SIGNAL mux_1053_nl : STD_LOGIC;
  SIGNAL mux_1050_nl : STD_LOGIC;
  SIGNAL or_1996_nl : STD_LOGIC;
  SIGNAL mux_1049_nl : STD_LOGIC;
  SIGNAL mux_1048_nl : STD_LOGIC;
  SIGNAL or_1994_nl : STD_LOGIC;
  SIGNAL mux_1047_nl : STD_LOGIC;
  SIGNAL mux_1046_nl : STD_LOGIC;
  SIGNAL mux_1045_nl : STD_LOGIC;
  SIGNAL mux_1043_nl : STD_LOGIC;
  SIGNAL mux_1042_nl : STD_LOGIC;
  SIGNAL mux_1072_nl : STD_LOGIC;
  SIGNAL mux_1071_nl : STD_LOGIC;
  SIGNAL mux_1070_nl : STD_LOGIC;
  SIGNAL nand_328_nl : STD_LOGIC;
  SIGNAL mux_1069_nl : STD_LOGIC;
  SIGNAL mux_1068_nl : STD_LOGIC;
  SIGNAL or_2016_nl : STD_LOGIC;
  SIGNAL or_2015_nl : STD_LOGIC;
  SIGNAL or_2014_nl : STD_LOGIC;
  SIGNAL mux_1067_nl : STD_LOGIC;
  SIGNAL mux_1066_nl : STD_LOGIC;
  SIGNAL or_2013_nl : STD_LOGIC;
  SIGNAL mux_1065_nl : STD_LOGIC;
  SIGNAL or_2008_nl : STD_LOGIC;
  SIGNAL mux_1064_nl : STD_LOGIC;
  SIGNAL or_2007_nl : STD_LOGIC;
  SIGNAL or_2006_nl : STD_LOGIC;
  SIGNAL nand_329_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_mux_22_nl : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_quantized_value_mux_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_mux_24_nl : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_quantized_value_mux_1_nl : STD_LOGIC_VECTOR (38
      DOWNTO 0);
  SIGNAL for_for_mux1h_5_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL for_for_for_for_nand_nl : STD_LOGIC;
  SIGNAL for_for_and_24_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_not_nl : STD_LOGIC;
  SIGNAL for_for_mux1h_6_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_attn_output_2D_not_3_nl : STD_LOGIC;
  SIGNAL mux_1099_nl : STD_LOGIC;
  SIGNAL mux_1097_nl : STD_LOGIC;
  SIGNAL mux_1095_nl : STD_LOGIC;
  SIGNAL or_2048_nl : STD_LOGIC;
  SIGNAL mux_1116_nl : STD_LOGIC;
  SIGNAL mux_1115_nl : STD_LOGIC;
  SIGNAL mux_1114_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_36_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_52_nl : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL for_for_and_22_nl : STD_LOGIC;
  SIGNAL mux_1119_nl : STD_LOGIC;
  SIGNAL mux_1118_nl : STD_LOGIC;
  SIGNAL mux_1117_nl : STD_LOGIC;
  SIGNAL or_2081_nl : STD_LOGIC;
  SIGNAL or_2080_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_28_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_nl : STD_LOGIC;
  SIGNAL and_521_nl : STD_LOGIC;
  SIGNAL and_523_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_29_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_1_nl : STD_LOGIC;
  SIGNAL and_527_nl : STD_LOGIC;
  SIGNAL and_529_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_31_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_3_nl : STD_LOGIC;
  SIGNAL and_531_nl : STD_LOGIC;
  SIGNAL and_533_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_33_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_5_nl : STD_LOGIC;
  SIGNAL and_535_nl : STD_LOGIC;
  SIGNAL and_537_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_and_35_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_7_nl : STD_LOGIC;
  SIGNAL and_539_nl : STD_LOGIC;
  SIGNAL and_541_nl : STD_LOGIC;
  SIGNAL mux_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL for_for_or_3_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL for_for_mux1h_13_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL for_for_or_4_nl : STD_LOGIC;
  SIGNAL for_for_and_28_nl : STD_LOGIC;
  SIGNAL or_nl : STD_LOGIC;
  SIGNAL nor_nl : STD_LOGIC;
  SIGNAL mux_1133_nl : STD_LOGIC;
  SIGNAL or_2087_nl : STD_LOGIC;
  SIGNAL mux1h_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL or_3215_nl : STD_LOGIC;
  SIGNAL not_4622_nl : STD_LOGIC;
  SIGNAL mux1h_1_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL or_3216_nl : STD_LOGIC;
  SIGNAL not_4624_nl : STD_LOGIC;
  SIGNAL mux1h_2_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL or_3217_nl : STD_LOGIC;
  SIGNAL not_4626_nl : STD_LOGIC;
  SIGNAL mux_1211_nl : STD_LOGIC;
  SIGNAL mux_1210_nl : STD_LOGIC;
  SIGNAL mux_1209_nl : STD_LOGIC;
  SIGNAL mux_1208_nl : STD_LOGIC;
  SIGNAL mux_1212_nl : STD_LOGIC;
  SIGNAL nor_1046_nl : STD_LOGIC;
  SIGNAL and_1597_nl : STD_LOGIC;
  SIGNAL mux_1235_nl : STD_LOGIC;
  SIGNAL mux_1234_nl : STD_LOGIC;
  SIGNAL mux_1233_nl : STD_LOGIC;
  SIGNAL mux_1232_nl : STD_LOGIC;
  SIGNAL mux_1231_nl : STD_LOGIC;
  SIGNAL mux_1230_nl : STD_LOGIC;
  SIGNAL mux_1228_nl : STD_LOGIC;
  SIGNAL mux_1227_nl : STD_LOGIC;
  SIGNAL mux_1226_nl : STD_LOGIC;
  SIGNAL mux_1225_nl : STD_LOGIC;
  SIGNAL mux_1224_nl : STD_LOGIC;
  SIGNAL mux_1223_nl : STD_LOGIC;
  SIGNAL or_2152_nl : STD_LOGIC;
  SIGNAL or_2151_nl : STD_LOGIC;
  SIGNAL or_2150_nl : STD_LOGIC;
  SIGNAL mux_1222_nl : STD_LOGIC;
  SIGNAL mux_1221_nl : STD_LOGIC;
  SIGNAL mux_1220_nl : STD_LOGIC;
  SIGNAL mux_1217_nl : STD_LOGIC;
  SIGNAL mux_1216_nl : STD_LOGIC;
  SIGNAL or_2145_nl : STD_LOGIC;
  SIGNAL mux_1215_nl : STD_LOGIC;
  SIGNAL mux_1214_nl : STD_LOGIC;
  SIGNAL mux_1213_nl : STD_LOGIC;
  SIGNAL or_2142_nl : STD_LOGIC;
  SIGNAL or_2140_nl : STD_LOGIC;
  SIGNAL or_2138_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_7_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_4_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_10_nl : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL mux_1310_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_proj_attention_2_1_16_16_4_4_q_proj_mux_12_nl
      : STD_LOGIC;
  SIGNAL mux_1308_nl : STD_LOGIC;
  SIGNAL or_3174_nl : STD_LOGIC;
  SIGNAL nand_344_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_and_2_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_i_mux1h_3_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_2_2_i_not_2_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_i_mux1h_6_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_and_10_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_38_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_10_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_39_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_11_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_40_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_12_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_41_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_13_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_42_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_14_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_43_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_15_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_44_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_16_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_1_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_1_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_24_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_17_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_18_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_26_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_19_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_27_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_20_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_28_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_21_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_29_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_22_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_30_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_23_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_2_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_2_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_10_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_24_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_11_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_25_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_12_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_26_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_13_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_27_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_14_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_28_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_15_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_29_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_16_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_30_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_3_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_3_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_17_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_31_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_18_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_32_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_19_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_33_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_20_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_34_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_21_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_35_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_22_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_36_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_23_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_37_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_4_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_4_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_31_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_38_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_32_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_39_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_33_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_40_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_34_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_41_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_35_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_42_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_36_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_43_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_37_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_44_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_5_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_5_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_45_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_45_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_46_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_46_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_47_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_47_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_48_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_48_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_49_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_49_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_50_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_50_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_51_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_51_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_6_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_6_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_52_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_52_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_53_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_53_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_54_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_54_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_55_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_55_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_56_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_56_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_57_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_57_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_58_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_58_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_7_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_7_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_59_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_59_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_60_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_60_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_61_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_61_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_62_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_62_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_63_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_63_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_64_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_64_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_65_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_65_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_8_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_8_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_66_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_66_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_67_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_67_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_68_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_68_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_69_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_69_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_70_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_70_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_71_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_71_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_72_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_72_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_9_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_9_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_73_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_73_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_74_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_74_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_75_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_75_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_76_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_76_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_77_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_77_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_78_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_78_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_79_nl : STD_LOGIC;
  SIGNAL INIT_2D_MEM_LOOP_2_mux_79_nl : STD_LOGIC;
  SIGNAL mux_1434_nl : STD_LOGIC;
  SIGNAL mux_1433_nl : STD_LOGIC;
  SIGNAL or_2335_nl : STD_LOGIC;
  SIGNAL mux_1432_nl : STD_LOGIC;
  SIGNAL mux_1431_nl : STD_LOGIC;
  SIGNAL mux_1430_nl : STD_LOGIC;
  SIGNAL mux_1429_nl : STD_LOGIC;
  SIGNAL mux_1428_nl : STD_LOGIC;
  SIGNAL nor_1105_nl : STD_LOGIC;
  SIGNAL or_2331_nl : STD_LOGIC;
  SIGNAL mux_1638_nl : STD_LOGIC;
  SIGNAL nand_71_nl : STD_LOGIC;
  SIGNAL or_2563_nl : STD_LOGIC;
  SIGNAL mux_1637_nl : STD_LOGIC;
  SIGNAL mux_1636_nl : STD_LOGIC;
  SIGNAL mux_1453_nl : STD_LOGIC;
  SIGNAL mux_1452_nl : STD_LOGIC;
  SIGNAL and_679_nl : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_3_nl : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_and_nl : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_4_nl : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_3_nl : STD_LOGIC;
  SIGNAL CACHE_UPDATE_LOOP_3_k_and_1_nl : STD_LOGIC;
  SIGNAL mux_1441_nl : STD_LOGIC;
  SIGNAL nor_1109_nl : STD_LOGIC;
  SIGNAL nor_1110_nl : STD_LOGIC;
  SIGNAL mux_1457_nl : STD_LOGIC;
  SIGNAL nor_1115_nl : STD_LOGIC;
  SIGNAL mux_1456_nl : STD_LOGIC;
  SIGNAL nand_350_nl : STD_LOGIC;
  SIGNAL or_2355_nl : STD_LOGIC;
  SIGNAL mux_1455_nl : STD_LOGIC;
  SIGNAL nor_1116_nl : STD_LOGIC;
  SIGNAL nor_1117_nl : STD_LOGIC;
  SIGNAL mux_1454_nl : STD_LOGIC;
  SIGNAL nor_1114_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_1_i_mux_1_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_and_36_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_mux1h_nl : STD_LOGIC;
  SIGNAL or_594_nl : STD_LOGIC;
  SIGNAL mux_1439_nl : STD_LOGIC;
  SIGNAL or_2342_nl : STD_LOGIC;
  SIGNAL mux_1438_nl : STD_LOGIC;
  SIGNAL nand_348_nl : STD_LOGIC;
  SIGNAL or_2341_nl : STD_LOGIC;
  SIGNAL mux_1437_nl : STD_LOGIC;
  SIGNAL or_2340_nl : STD_LOGIC;
  SIGNAL or_2339_nl : STD_LOGIC;
  SIGNAL mux_1490_nl : STD_LOGIC;
  SIGNAL nand_126_nl : STD_LOGIC;
  SIGNAL and_688_nl : STD_LOGIC;
  SIGNAL and_693_nl : STD_LOGIC;
  SIGNAL and_704_nl : STD_LOGIC;
  SIGNAL and_709_nl : STD_LOGIC;
  SIGNAL and_713_nl : STD_LOGIC;
  SIGNAL and_717_nl : STD_LOGIC;
  SIGNAL and_721_nl : STD_LOGIC;
  SIGNAL and_725_nl : STD_LOGIC;
  SIGNAL and_729_nl : STD_LOGIC;
  SIGNAL and_733_nl : STD_LOGIC;
  SIGNAL and_737_nl : STD_LOGIC;
  SIGNAL and_741_nl : STD_LOGIC;
  SIGNAL and_749_nl : STD_LOGIC;
  SIGNAL and_753_nl : STD_LOGIC;
  SIGNAL or_2443_nl : STD_LOGIC;
  SIGNAL mux_1498_nl : STD_LOGIC;
  SIGNAL mux_1497_nl : STD_LOGIC;
  SIGNAL or_2429_nl : STD_LOGIC;
  SIGNAL mux_1496_nl : STD_LOGIC;
  SIGNAL or_2426_nl : STD_LOGIC;
  SIGNAL mux_1495_nl : STD_LOGIC;
  SIGNAL mux_1494_nl : STD_LOGIC;
  SIGNAL mux_1493_nl : STD_LOGIC;
  SIGNAL mux_1492_nl : STD_LOGIC;
  SIGNAL nand_354_nl : STD_LOGIC;
  SIGNAL nand_355_nl : STD_LOGIC;
  SIGNAL mux_1511_nl : STD_LOGIC;
  SIGNAL mux_1510_nl : STD_LOGIC;
  SIGNAL or_2442_nl : STD_LOGIC;
  SIGNAL mux_1509_nl : STD_LOGIC;
  SIGNAL mux_1508_nl : STD_LOGIC;
  SIGNAL mux_1507_nl : STD_LOGIC;
  SIGNAL or_2441_nl : STD_LOGIC;
  SIGNAL mux_1505_nl : STD_LOGIC;
  SIGNAL or_2438_nl : STD_LOGIC;
  SIGNAL nand_64_nl : STD_LOGIC;
  SIGNAL mux_1504_nl : STD_LOGIC;
  SIGNAL mux_1503_nl : STD_LOGIC;
  SIGNAL or_2436_nl : STD_LOGIC;
  SIGNAL nand_63_nl : STD_LOGIC;
  SIGNAL mux_1502_nl : STD_LOGIC;
  SIGNAL mux_1501_nl : STD_LOGIC;
  SIGNAL mux_1500_nl : STD_LOGIC;
  SIGNAL or_2431_nl : STD_LOGIC;
  SIGNAL mux_1533_nl : STD_LOGIC;
  SIGNAL mux_1532_nl : STD_LOGIC;
  SIGNAL mux_1531_nl : STD_LOGIC;
  SIGNAL mux_1530_nl : STD_LOGIC;
  SIGNAL mux_1529_nl : STD_LOGIC;
  SIGNAL or_2459_nl : STD_LOGIC;
  SIGNAL mux_1528_nl : STD_LOGIC;
  SIGNAL mux_1527_nl : STD_LOGIC;
  SIGNAL or_2458_nl : STD_LOGIC;
  SIGNAL mux_1526_nl : STD_LOGIC;
  SIGNAL mux_1525_nl : STD_LOGIC;
  SIGNAL mux_1524_nl : STD_LOGIC;
  SIGNAL mux_1523_nl : STD_LOGIC;
  SIGNAL mux_1521_nl : STD_LOGIC;
  SIGNAL mux_1520_nl : STD_LOGIC;
  SIGNAL mux_1518_nl : STD_LOGIC;
  SIGNAL mux_1517_nl : STD_LOGIC;
  SIGNAL or_2448_nl : STD_LOGIC;
  SIGNAL or_2446_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_1_i_mux1h_5_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_and_1_nl : STD_LOGIC;
  SIGNAL and_755_nl : STD_LOGIC;
  SIGNAL nor_1136_nl : STD_LOGIC;
  SIGNAL mux_1491_nl : STD_LOGIC;
  SIGNAL nand_353_nl : STD_LOGIC;
  SIGNAL and_757_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_1_i_or_nl : STD_LOGIC;
  SIGNAL mux_1516_nl : STD_LOGIC;
  SIGNAL nand_356_nl : STD_LOGIC;
  SIGNAL mux_1515_nl : STD_LOGIC;
  SIGNAL mux_1514_nl : STD_LOGIC;
  SIGNAL mux_1537_nl : STD_LOGIC;
  SIGNAL mux_1536_nl : STD_LOGIC;
  SIGNAL nor_1141_nl : STD_LOGIC;
  SIGNAL nor_1142_nl : STD_LOGIC;
  SIGNAL nor_1143_nl : STD_LOGIC;
  SIGNAL mux_1534_nl : STD_LOGIC;
  SIGNAL or_2463_nl : STD_LOGIC;
  SIGNAL or_2461_nl : STD_LOGIC;
  SIGNAL mux_1541_nl : STD_LOGIC;
  SIGNAL mux_1540_nl : STD_LOGIC;
  SIGNAL mux_1539_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_4_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4557_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_8_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4558_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_12_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4559_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_16_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4560_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_20_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4561_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_21_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4562_nl : STD_LOGIC;
  SIGNAL mux_1554_nl : STD_LOGIC;
  SIGNAL and_1652_nl : STD_LOGIC;
  SIGNAL mux_1552_nl : STD_LOGIC;
  SIGNAL mux_1550_nl : STD_LOGIC;
  SIGNAL or_2479_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_5_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_779_nl : STD_LOGIC;
  SIGNAL mux_1561_nl : STD_LOGIC;
  SIGNAL mux_1560_nl : STD_LOGIC;
  SIGNAL mux_1558_nl : STD_LOGIC;
  SIGNAL mux_1556_nl : STD_LOGIC;
  SIGNAL and_1653_nl : STD_LOGIC;
  SIGNAL and_783_nl : STD_LOGIC;
  SIGNAL and_790_nl : STD_LOGIC;
  SIGNAL not_4472_nl : STD_LOGIC;
  SIGNAL mux_1564_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_35_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4441_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_34_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4440_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_33_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4439_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_32_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4438_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_31_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4437_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_30_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4436_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_29_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4435_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_28_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4434_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_27_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4433_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_26_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4432_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_25_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4431_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_24_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4430_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_23_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4429_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_22_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4428_nl : STD_LOGIC;
  SIGNAL mux_1581_nl : STD_LOGIC;
  SIGNAL or_2494_nl : STD_LOGIC;
  SIGNAL mux_1580_nl : STD_LOGIC;
  SIGNAL or_2493_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_21_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4427_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_20_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4426_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_19_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4425_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_18_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4424_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_40_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4423_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_17_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4422_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_42_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4421_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_43_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4420_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_44_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4419_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_45_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4418_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_46_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4417_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_47_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4416_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_16_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4415_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_l_GEMM_3D_FLOAT_LOOP_4_l_mux_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_l_mux1h_13_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_or_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_mux_23_nl : STD_LOGIC;
  SIGNAL and_1254_nl : STD_LOGIC;
  SIGNAL mux_2245_nl : STD_LOGIC;
  SIGNAL mux_2244_nl : STD_LOGIC;
  SIGNAL mux_2243_nl : STD_LOGIC;
  SIGNAL mux_2242_nl : STD_LOGIC;
  SIGNAL and_1810_nl : STD_LOGIC;
  SIGNAL mux_2241_nl : STD_LOGIC;
  SIGNAL nor_1320_nl : STD_LOGIC;
  SIGNAL mux_2240_nl : STD_LOGIC;
  SIGNAL nor_1316_nl : STD_LOGIC;
  SIGNAL mux_2239_nl : STD_LOGIC;
  SIGNAL and_1809_nl : STD_LOGIC;
  SIGNAL nor_1321_nl : STD_LOGIC;
  SIGNAL mux_2238_nl : STD_LOGIC;
  SIGNAL or_3033_nl : STD_LOGIC;
  SIGNAL or_3032_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_l_or_1_nl : STD_LOGIC;
  SIGNAL or_2566_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_26_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_939_nl : STD_LOGIC;
  SIGNAL not_4471_nl : STD_LOGIC;
  SIGNAL mux_1641_nl : STD_LOGIC;
  SIGNAL or_3192_nl : STD_LOGIC;
  SIGNAL mux_1640_nl : STD_LOGIC;
  SIGNAL or_3191_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_28_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_941_nl : STD_LOGIC;
  SIGNAL not_4470_nl : STD_LOGIC;
  SIGNAL mux_1644_nl : STD_LOGIC;
  SIGNAL or_3195_nl : STD_LOGIC;
  SIGNAL mux_1643_nl : STD_LOGIC;
  SIGNAL or_3194_nl : STD_LOGIC;
  SIGNAL or_2576_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_30_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_943_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_nand_nl : STD_LOGIC;
  SIGNAL mux_1660_nl : STD_LOGIC;
  SIGNAL mux_1659_nl : STD_LOGIC;
  SIGNAL mux_1657_nl : STD_LOGIC;
  SIGNAL mux_1655_nl : STD_LOGIC;
  SIGNAL nor_466_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_and_81_nl : STD_LOGIC;
  SIGNAL and_945_nl : STD_LOGIC;
  SIGNAL not_4469_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_32_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_946_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_nand_2_nl : STD_LOGIC;
  SIGNAL mux_1676_nl : STD_LOGIC;
  SIGNAL mux_1675_nl : STD_LOGIC;
  SIGNAL mux_1673_nl : STD_LOGIC;
  SIGNAL mux_1671_nl : STD_LOGIC;
  SIGNAL and_1684_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_and_83_nl : STD_LOGIC;
  SIGNAL and_948_nl : STD_LOGIC;
  SIGNAL not_4468_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_34_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_949_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_nand_4_nl : STD_LOGIC;
  SIGNAL mux_1692_nl : STD_LOGIC;
  SIGNAL mux_1691_nl : STD_LOGIC;
  SIGNAL mux_1689_nl : STD_LOGIC;
  SIGNAL mux_1687_nl : STD_LOGIC;
  SIGNAL or_2589_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_and_85_nl : STD_LOGIC;
  SIGNAL and_951_nl : STD_LOGIC;
  SIGNAL not_4467_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_36_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_952_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_nand_6_nl : STD_LOGIC;
  SIGNAL mux_1708_nl : STD_LOGIC;
  SIGNAL mux_1707_nl : STD_LOGIC;
  SIGNAL mux_1705_nl : STD_LOGIC;
  SIGNAL mux_1703_nl : STD_LOGIC;
  SIGNAL nand_367_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_and_87_nl : STD_LOGIC;
  SIGNAL and_954_nl : STD_LOGIC;
  SIGNAL not_4466_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_38_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_955_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_nand_8_nl : STD_LOGIC;
  SIGNAL mux_1724_nl : STD_LOGIC;
  SIGNAL mux_1723_nl : STD_LOGIC;
  SIGNAL mux_1721_nl : STD_LOGIC;
  SIGNAL mux_1719_nl : STD_LOGIC;
  SIGNAL and_1697_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_and_89_nl : STD_LOGIC;
  SIGNAL and_957_nl : STD_LOGIC;
  SIGNAL not_4465_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_40_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_958_nl : STD_LOGIC;
  SIGNAL not_4464_nl : STD_LOGIC;
  SIGNAL mux_1727_nl : STD_LOGIC;
  SIGNAL or_3197_nl : STD_LOGIC;
  SIGNAL mux_1726_nl : STD_LOGIC;
  SIGNAL nand_81_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_42_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_960_nl : STD_LOGIC;
  SIGNAL mux_1743_nl : STD_LOGIC;
  SIGNAL mux_1742_nl : STD_LOGIC;
  SIGNAL mux_1740_nl : STD_LOGIC;
  SIGNAL mux_1738_nl : STD_LOGIC;
  SIGNAL or_2611_nl : STD_LOGIC;
  SIGNAL and_962_nl : STD_LOGIC;
  SIGNAL not_4463_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_44_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_963_nl : STD_LOGIC;
  SIGNAL mux_1759_nl : STD_LOGIC;
  SIGNAL mux_1758_nl : STD_LOGIC;
  SIGNAL mux_1756_nl : STD_LOGIC;
  SIGNAL mux_1754_nl : STD_LOGIC;
  SIGNAL or_2617_nl : STD_LOGIC;
  SIGNAL and_965_nl : STD_LOGIC;
  SIGNAL not_4462_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_46_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_966_nl : STD_LOGIC;
  SIGNAL mux_1775_nl : STD_LOGIC;
  SIGNAL mux_1774_nl : STD_LOGIC;
  SIGNAL mux_1772_nl : STD_LOGIC;
  SIGNAL mux_1770_nl : STD_LOGIC;
  SIGNAL nor_500_nl : STD_LOGIC;
  SIGNAL and_968_nl : STD_LOGIC;
  SIGNAL not_4461_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_48_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_969_nl : STD_LOGIC;
  SIGNAL mux_1791_nl : STD_LOGIC;
  SIGNAL mux_1790_nl : STD_LOGIC;
  SIGNAL mux_1788_nl : STD_LOGIC;
  SIGNAL mux_1786_nl : STD_LOGIC;
  SIGNAL or_2492_nl : STD_LOGIC;
  SIGNAL and_971_nl : STD_LOGIC;
  SIGNAL not_4460_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_50_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_972_nl : STD_LOGIC;
  SIGNAL mux_1807_nl : STD_LOGIC;
  SIGNAL mux_1806_nl : STD_LOGIC;
  SIGNAL mux_1804_nl : STD_LOGIC;
  SIGNAL mux_1802_nl : STD_LOGIC;
  SIGNAL or_2497_nl : STD_LOGIC;
  SIGNAL and_974_nl : STD_LOGIC;
  SIGNAL not_4459_nl : STD_LOGIC;
  SIGNAL mux_1811_nl : STD_LOGIC;
  SIGNAL mux_1810_nl : STD_LOGIC;
  SIGNAL or_2638_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_43_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4458_nl : STD_LOGIC;
  SIGNAL mux_1816_nl : STD_LOGIC;
  SIGNAL mux_1815_nl : STD_LOGIC;
  SIGNAL mux_1814_nl : STD_LOGIC;
  SIGNAL mux_1813_nl : STD_LOGIC;
  SIGNAL or_2491_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_42_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4457_nl : STD_LOGIC;
  SIGNAL mux_1825_nl : STD_LOGIC;
  SIGNAL mux_1824_nl : STD_LOGIC;
  SIGNAL mux_1823_nl : STD_LOGIC;
  SIGNAL mux_1822_nl : STD_LOGIC;
  SIGNAL or_2490_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_41_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4456_nl : STD_LOGIC;
  SIGNAL mux_1834_nl : STD_LOGIC;
  SIGNAL mux_1833_nl : STD_LOGIC;
  SIGNAL mux_1832_nl : STD_LOGIC;
  SIGNAL mux_1831_nl : STD_LOGIC;
  SIGNAL nor_514_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_40_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4455_nl : STD_LOGIC;
  SIGNAL mux_1843_nl : STD_LOGIC;
  SIGNAL mux_1842_nl : STD_LOGIC;
  SIGNAL mux_1841_nl : STD_LOGIC;
  SIGNAL mux_1840_nl : STD_LOGIC;
  SIGNAL and_1727_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_39_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4454_nl : STD_LOGIC;
  SIGNAL mux_1852_nl : STD_LOGIC;
  SIGNAL mux_1851_nl : STD_LOGIC;
  SIGNAL mux_1850_nl : STD_LOGIC;
  SIGNAL mux_1849_nl : STD_LOGIC;
  SIGNAL or_2653_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_38_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4453_nl : STD_LOGIC;
  SIGNAL mux_1861_nl : STD_LOGIC;
  SIGNAL mux_1860_nl : STD_LOGIC;
  SIGNAL mux_1859_nl : STD_LOGIC;
  SIGNAL mux_1858_nl : STD_LOGIC;
  SIGNAL nand_369_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_37_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4452_nl : STD_LOGIC;
  SIGNAL mux_1870_nl : STD_LOGIC;
  SIGNAL mux_1869_nl : STD_LOGIC;
  SIGNAL mux_1868_nl : STD_LOGIC;
  SIGNAL mux_1867_nl : STD_LOGIC;
  SIGNAL and_1658_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_36_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4451_nl : STD_LOGIC;
  SIGNAL mux_1878_nl : STD_LOGIC;
  SIGNAL mux_1877_nl : STD_LOGIC;
  SIGNAL mux_1876_nl : STD_LOGIC;
  SIGNAL mux_1875_nl : STD_LOGIC;
  SIGNAL mux_1874_nl : STD_LOGIC;
  SIGNAL and_1733_nl : STD_LOGIC;
  SIGNAL mux_1873_nl : STD_LOGIC;
  SIGNAL or_2664_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_35_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4450_nl : STD_LOGIC;
  SIGNAL mux_1887_nl : STD_LOGIC;
  SIGNAL mux_1886_nl : STD_LOGIC;
  SIGNAL mux_1885_nl : STD_LOGIC;
  SIGNAL mux_1884_nl : STD_LOGIC;
  SIGNAL nor_524_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_34_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4449_nl : STD_LOGIC;
  SIGNAL mux_1896_nl : STD_LOGIC;
  SIGNAL mux_1895_nl : STD_LOGIC;
  SIGNAL mux_1894_nl : STD_LOGIC;
  SIGNAL mux_1893_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_33_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4448_nl : STD_LOGIC;
  SIGNAL mux_1905_nl : STD_LOGIC;
  SIGNAL mux_1904_nl : STD_LOGIC;
  SIGNAL mux_1903_nl : STD_LOGIC;
  SIGNAL mux_1902_nl : STD_LOGIC;
  SIGNAL or_2675_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_32_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4447_nl : STD_LOGIC;
  SIGNAL mux_1914_nl : STD_LOGIC;
  SIGNAL mux_1913_nl : STD_LOGIC;
  SIGNAL mux_1912_nl : STD_LOGIC;
  SIGNAL mux_1911_nl : STD_LOGIC;
  SIGNAL nor_441_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_31_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4446_nl : STD_LOGIC;
  SIGNAL mux_1923_nl : STD_LOGIC;
  SIGNAL mux_1922_nl : STD_LOGIC;
  SIGNAL mux_1921_nl : STD_LOGIC;
  SIGNAL mux_1920_nl : STD_LOGIC;
  SIGNAL and_1656_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_30_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4445_nl : STD_LOGIC;
  SIGNAL mux_1932_nl : STD_LOGIC;
  SIGNAL mux_1931_nl : STD_LOGIC;
  SIGNAL mux_1930_nl : STD_LOGIC;
  SIGNAL mux_1929_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_29_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4444_nl : STD_LOGIC;
  SIGNAL mux_1941_nl : STD_LOGIC;
  SIGNAL mux_1940_nl : STD_LOGIC;
  SIGNAL mux_1939_nl : STD_LOGIC;
  SIGNAL mux_1938_nl : STD_LOGIC;
  SIGNAL or_2487_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_66_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_1025_nl : STD_LOGIC;
  SIGNAL not_4563_nl : STD_LOGIC;
  SIGNAL mux_1946_nl : STD_LOGIC;
  SIGNAL nor_533_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_67_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_1031_nl : STD_LOGIC;
  SIGNAL not_4564_nl : STD_LOGIC;
  SIGNAL mux_1947_nl : STD_LOGIC;
  SIGNAL nor_535_nl : STD_LOGIC;
  SIGNAL mux_1965_nl : STD_LOGIC;
  SIGNAL mux_1964_nl : STD_LOGIC;
  SIGNAL mux_1962_nl : STD_LOGIC;
  SIGNAL mux_1961_nl : STD_LOGIC;
  SIGNAL mux_1960_nl : STD_LOGIC;
  SIGNAL mux_1959_nl : STD_LOGIC;
  SIGNAL mux_1958_nl : STD_LOGIC;
  SIGNAL mux_1957_nl : STD_LOGIC;
  SIGNAL mux_1954_nl : STD_LOGIC;
  SIGNAL nor_540_nl : STD_LOGIC;
  SIGNAL mux_1950_nl : STD_LOGIC;
  SIGNAL or_2696_nl : STD_LOGIC;
  SIGNAL mux_1949_nl : STD_LOGIC;
  SIGNAL mux_1948_nl : STD_LOGIC;
  SIGNAL or_2695_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_68_nl : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_118_nl : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL not_4443_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_69_nl : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_119_nl : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL not_4565_nl : STD_LOGIC;
  SIGNAL mux_1973_nl : STD_LOGIC;
  SIGNAL mux_1972_nl : STD_LOGIC;
  SIGNAL and_1753_nl : STD_LOGIC;
  SIGNAL mux_1971_nl : STD_LOGIC;
  SIGNAL mux_1970_nl : STD_LOGIC;
  SIGNAL nor_1203_nl : STD_LOGIC;
  SIGNAL nor_1204_nl : STD_LOGIC;
  SIGNAL and_1749_nl : STD_LOGIC;
  SIGNAL mux_1969_nl : STD_LOGIC;
  SIGNAL nor_1201_nl : STD_LOGIC;
  SIGNAL nor_1202_nl : STD_LOGIC;
  SIGNAL nor_1206_nl : STD_LOGIC;
  SIGNAL mux_1968_nl : STD_LOGIC;
  SIGNAL mux_1967_nl : STD_LOGIC;
  SIGNAL and_1754_nl : STD_LOGIC;
  SIGNAL nor_1208_nl : STD_LOGIC;
  SIGNAL mux_1985_nl : STD_LOGIC;
  SIGNAL mux_1984_nl : STD_LOGIC;
  SIGNAL mux_1983_nl : STD_LOGIC;
  SIGNAL mux_1982_nl : STD_LOGIC;
  SIGNAL nor_551_nl : STD_LOGIC;
  SIGNAL mux_1978_nl : STD_LOGIC;
  SIGNAL mux_1977_nl : STD_LOGIC;
  SIGNAL mux_1976_nl : STD_LOGIC;
  SIGNAL or_2712_nl : STD_LOGIC;
  SIGNAL mux_1975_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_70_nl : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL not_5074_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_128_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_129_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_130_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_131_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_132_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_133_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_134_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_135_nl : STD_LOGIC;
  SIGNAL mux_1998_nl : STD_LOGIC;
  SIGNAL mux_1997_nl : STD_LOGIC;
  SIGNAL mux_1996_nl : STD_LOGIC;
  SIGNAL mux_1995_nl : STD_LOGIC;
  SIGNAL mux_1994_nl : STD_LOGIC;
  SIGNAL nor_552_nl : STD_LOGIC;
  SIGNAL mux_1992_nl : STD_LOGIC;
  SIGNAL mux_1991_nl : STD_LOGIC;
  SIGNAL mux_1989_nl : STD_LOGIC;
  SIGNAL mux_1988_nl : STD_LOGIC;
  SIGNAL or_2716_nl : STD_LOGIC;
  SIGNAL mux_1987_nl : STD_LOGIC;
  SIGNAL or_2715_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_71_nl : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL not_5066_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_120_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_121_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_122_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_123_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_124_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_125_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_126_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_127_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_72_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4566_nl : STD_LOGIC;
  SIGNAL mux_2012_nl : STD_LOGIC;
  SIGNAL mux_2011_nl : STD_LOGIC;
  SIGNAL nand_93_nl : STD_LOGIC;
  SIGNAL mux_2010_nl : STD_LOGIC;
  SIGNAL mux_2009_nl : STD_LOGIC;
  SIGNAL mux_2008_nl : STD_LOGIC;
  SIGNAL mux_2007_nl : STD_LOGIC;
  SIGNAL nand_92_nl : STD_LOGIC;
  SIGNAL mux_2006_nl : STD_LOGIC;
  SIGNAL mux_2005_nl : STD_LOGIC;
  SIGNAL mux_2003_nl : STD_LOGIC;
  SIGNAL mux_2002_nl : STD_LOGIC;
  SIGNAL and_1759_nl : STD_LOGIC;
  SIGNAL mux_2001_nl : STD_LOGIC;
  SIGNAL mux_2000_nl : STD_LOGIC;
  SIGNAL or_2720_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_73_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4567_nl : STD_LOGIC;
  SIGNAL mux_2022_nl : STD_LOGIC;
  SIGNAL mux_2021_nl : STD_LOGIC;
  SIGNAL mux_2020_nl : STD_LOGIC;
  SIGNAL mux_2019_nl : STD_LOGIC;
  SIGNAL mux_2018_nl : STD_LOGIC;
  SIGNAL or_2733_nl : STD_LOGIC;
  SIGNAL and_1763_nl : STD_LOGIC;
  SIGNAL mux_2017_nl : STD_LOGIC;
  SIGNAL mux_2016_nl : STD_LOGIC;
  SIGNAL mux_2033_nl : STD_LOGIC;
  SIGNAL mux_2031_nl : STD_LOGIC;
  SIGNAL mux_2030_nl : STD_LOGIC;
  SIGNAL mux_2029_nl : STD_LOGIC;
  SIGNAL mux_2028_nl : STD_LOGIC;
  SIGNAL or_2741_nl : STD_LOGIC;
  SIGNAL mux_2027_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_74_nl : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL not_5054_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_117_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_67_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_152_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_88_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_153_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_89_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_154_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_90_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_155_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_91_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_156_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_92_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_157_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_93_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_158_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_94_nl : STD_LOGIC;
  SIGNAL mux_2036_nl : STD_LOGIC;
  SIGNAL nor_410_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_75_nl : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL not_4569_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_116_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_144_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_145_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_146_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_147_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_148_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_149_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_150_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_151_nl : STD_LOGIC;
  SIGNAL not_5062_nl : STD_LOGIC;
  SIGNAL mux_2037_nl : STD_LOGIC;
  SIGNAL and_1626_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_76_nl : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL not_5088_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_136_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_137_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_138_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_139_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_140_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_141_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_142_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_143_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_77_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_1064_nl : STD_LOGIC;
  SIGNAL not_4571_nl : STD_LOGIC;
  SIGNAL mux_2038_nl : STD_LOGIC;
  SIGNAL nor_796_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_78_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_1066_nl : STD_LOGIC;
  SIGNAL not_4572_nl : STD_LOGIC;
  SIGNAL mux_2039_nl : STD_LOGIC;
  SIGNAL and_1420_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_79_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_1068_nl : STD_LOGIC;
  SIGNAL not_4573_nl : STD_LOGIC;
  SIGNAL mux_2040_nl : STD_LOGIC;
  SIGNAL and_1613_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_80_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_1071_nl : STD_LOGIC;
  SIGNAL and_1074_nl : STD_LOGIC;
  SIGNAL not_4574_nl : STD_LOGIC;
  SIGNAL mux_2051_nl : STD_LOGIC;
  SIGNAL mux_2049_nl : STD_LOGIC;
  SIGNAL mux_2048_nl : STD_LOGIC;
  SIGNAL mux_2047_nl : STD_LOGIC;
  SIGNAL mux_2046_nl : STD_LOGIC;
  SIGNAL or_2751_nl : STD_LOGIC;
  SIGNAL mux_2045_nl : STD_LOGIC;
  SIGNAL and_1660_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_81_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_1075_nl : STD_LOGIC;
  SIGNAL not_4575_nl : STD_LOGIC;
  SIGNAL mux_2052_nl : STD_LOGIC;
  SIGNAL or_2753_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_82_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_1081_nl : STD_LOGIC;
  SIGNAL not_4576_nl : STD_LOGIC;
  SIGNAL mux_2053_nl : STD_LOGIC;
  SIGNAL or_2281_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_83_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_1083_nl : STD_LOGIC;
  SIGNAL not_4577_nl : STD_LOGIC;
  SIGNAL mux_2054_nl : STD_LOGIC;
  SIGNAL or_2292_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux1h_84_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL and_1086_nl : STD_LOGIC;
  SIGNAL not_4578_nl : STD_LOGIC;
  SIGNAL mux_2055_nl : STD_LOGIC;
  SIGNAL or_2756_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_51_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL and_1089_nl : STD_LOGIC;
  SIGNAL mux_2056_nl : STD_LOGIC;
  SIGNAL or_2757_nl : STD_LOGIC;
  SIGNAL not_4414_nl : STD_LOGIC;
  SIGNAL mux_2059_nl : STD_LOGIC;
  SIGNAL or_3200_nl : STD_LOGIC;
  SIGNAL mux_2058_nl : STD_LOGIC;
  SIGNAL and_1090_nl : STD_LOGIC;
  SIGNAL mux_2057_nl : STD_LOGIC;
  SIGNAL nor_1217_nl : STD_LOGIC;
  SIGNAL or_3201_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_52_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4413_nl : STD_LOGIC;
  SIGNAL mux_2063_nl : STD_LOGIC;
  SIGNAL or_2764_nl : STD_LOGIC;
  SIGNAL mux_2062_nl : STD_LOGIC;
  SIGNAL or_2763_nl : STD_LOGIC;
  SIGNAL mux_2061_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_53_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL and_1097_nl : STD_LOGIC;
  SIGNAL mux_2064_nl : STD_LOGIC;
  SIGNAL or_2765_nl : STD_LOGIC;
  SIGNAL not_4412_nl : STD_LOGIC;
  SIGNAL mux_2068_nl : STD_LOGIC;
  SIGNAL mux_2065_nl : STD_LOGIC;
  SIGNAL nand_370_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_54_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_55_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4579_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_56_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_36_nl : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL not_4580_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_57_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_mux_33_nl : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_38_nl : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL not_4581_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_58_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_39_nl : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL not_4582_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_59_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4583_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_60_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4584_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_61_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4585_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_62_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4586_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_63_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4587_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux1h_64_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4588_nl : STD_LOGIC;
  SIGNAL mux_2088_nl : STD_LOGIC;
  SIGNAL mux_2087_nl : STD_LOGIC;
  SIGNAL mux_2086_nl : STD_LOGIC;
  SIGNAL mux_1542_nl : STD_LOGIC;
  SIGNAL nand_357_nl : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_nl
      : STD_LOGIC;
  SIGNAL mux_2099_nl : STD_LOGIC;
  SIGNAL mux_2098_nl : STD_LOGIC;
  SIGNAL or_2799_nl : STD_LOGIC;
  SIGNAL mux_2097_nl : STD_LOGIC;
  SIGNAL mux_2096_nl : STD_LOGIC;
  SIGNAL mux_2095_nl : STD_LOGIC;
  SIGNAL mux_2094_nl : STD_LOGIC;
  SIGNAL mux_2093_nl : STD_LOGIC;
  SIGNAL mux_2091_nl : STD_LOGIC;
  SIGNAL mux_2090_nl : STD_LOGIC;
  SIGNAL or_2787_nl : STD_LOGIC;
  SIGNAL or_2786_nl : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_1_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_APPLY_ROTARY_POS_EMB_LOOP_3_nor_nl : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_or_2_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_66_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_74_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_75_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_76_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_77_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_78_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_79_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_80_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_61_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_81_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_82_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_83_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_84_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_85_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_86_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_87_nl : STD_LOGIC;
  SIGNAL mux_2102_nl : STD_LOGIC;
  SIGNAL nand_283_nl : STD_LOGIC;
  SIGNAL mux_2104_nl : STD_LOGIC;
  SIGNAL mux_2103_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_32_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_70_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_71_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_72_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_50_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_51_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_52_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_53_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_54_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_55_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_56_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_57_nl : STD_LOGIC;
  SIGNAL mux_2108_nl : STD_LOGIC;
  SIGNAL nand_285_nl : STD_LOGIC;
  SIGNAL or_3153_nl : STD_LOGIC;
  SIGNAL mux_2107_nl : STD_LOGIC;
  SIGNAL or_2828_nl : STD_LOGIC;
  SIGNAL and_1184_nl : STD_LOGIC;
  SIGNAL mux_2109_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_1_mux_4_nl : STD_LOGIC;
  SIGNAL mux_2127_nl : STD_LOGIC;
  SIGNAL mux_2126_nl : STD_LOGIC;
  SIGNAL mux_2125_nl : STD_LOGIC;
  SIGNAL mux_2124_nl : STD_LOGIC;
  SIGNAL mux_2123_nl : STD_LOGIC;
  SIGNAL mux_2122_nl : STD_LOGIC;
  SIGNAL mux_2120_nl : STD_LOGIC;
  SIGNAL mux_2114_nl : STD_LOGIC;
  SIGNAL or_2840_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_and_7_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_and_5_nl : STD_LOGIC;
  SIGNAL mux_2128_nl : STD_LOGIC;
  SIGNAL mux_2130_nl : STD_LOGIC;
  SIGNAL mux_2129_nl : STD_LOGIC;
  SIGNAL mux_2131_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_mux1h_40_nl : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_or_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_33_nl : STD_LOGIC;
  SIGNAL not_4510_nl : STD_LOGIC;
  SIGNAL mux_2156_nl : STD_LOGIC;
  SIGNAL mux_2155_nl : STD_LOGIC;
  SIGNAL nor_1240_nl : STD_LOGIC;
  SIGNAL nor_1241_nl : STD_LOGIC;
  SIGNAL nor_1242_nl : STD_LOGIC;
  SIGNAL mux_2154_nl : STD_LOGIC;
  SIGNAL nor_1243_nl : STD_LOGIC;
  SIGNAL nor_1244_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_mux1h_41_nl : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL not_4483_nl : STD_LOGIC;
  SIGNAL mux_2159_nl : STD_LOGIC;
  SIGNAL mux_2158_nl : STD_LOGIC;
  SIGNAL nor_1245_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_mux1h_42_nl : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL not_4482_nl : STD_LOGIC;
  SIGNAL mux_2182_nl : STD_LOGIC;
  SIGNAL mux_2181_nl : STD_LOGIC;
  SIGNAL nor_1256_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_mux1h_43_nl : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_or_5_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_35_nl : STD_LOGIC;
  SIGNAL not_4511_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_mux1h_44_nl : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL not_4512_nl : STD_LOGIC;
  SIGNAL mux_2198_nl : STD_LOGIC;
  SIGNAL mux_2197_nl : STD_LOGIC;
  SIGNAL nor_1272_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_mux1h_45_nl : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL not_4513_nl : STD_LOGIC;
  SIGNAL mux_2204_nl : STD_LOGIC;
  SIGNAL mux_2203_nl : STD_LOGIC;
  SIGNAL nor_1283_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_mux1h_46_nl : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL not_4514_nl : STD_LOGIC;
  SIGNAL mux_2210_nl : STD_LOGIC;
  SIGNAL mux_2209_nl : STD_LOGIC;
  SIGNAL nor_1294_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_mux1h_47_nl : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_q_embed_or_6_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_and_37_nl : STD_LOGIC;
  SIGNAL not_4515_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_q_embed_mux1h_48_nl : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL not_4516_nl : STD_LOGIC;
  SIGNAL mux_2226_nl : STD_LOGIC;
  SIGNAL mux_2225_nl : STD_LOGIC;
  SIGNAL nor_1310_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_95_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_96_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_APPLY_ROTARY_POS_EMB_LOOP_6_or_7_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_97_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_98_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_99_nl : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_100_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux_101_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_35_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_not_28_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_34_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_not_27_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_33_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_not_26_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_32_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_not_25_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_31_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_not_24_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_30_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_not_23_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_29_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_not_22_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_28_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_not_21_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_27_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_not_20_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_26_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_not_19_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_25_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_not_18_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_3_and_24_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_3_not_17_nl : STD_LOGIC;
  SIGNAL mux_2237_nl : STD_LOGIC;
  SIGNAL mux_1543_nl : STD_LOGIC;
  SIGNAL mux_2248_nl : STD_LOGIC;
  SIGNAL nor_1319_nl : STD_LOGIC;
  SIGNAL mux_2250_nl : STD_LOGIC;
  SIGNAL mux_2249_nl : STD_LOGIC;
  SIGNAL mux_2258_nl : STD_LOGIC;
  SIGNAL mux_2257_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_nl : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL not_4589_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_44_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4590_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_36_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4591_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_45_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4592_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_37_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4593_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_46_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4594_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_38_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4595_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_47_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4596_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_39_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4597_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_48_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4598_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_40_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4599_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_49_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4600_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_41_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4601_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_50_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4602_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_42_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4603_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_51_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4604_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_43_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4605_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_52_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4606_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_44_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4607_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_53_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4608_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_45_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4609_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_54_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4610_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_46_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4611_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_55_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4612_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_47_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4613_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_56_nl : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL not_5055_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_60_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_61_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_62_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_63_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_64_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_65_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_66_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_67_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_48_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4615_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_57_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4616_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_49_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4617_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_58_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4618_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_proj_re_mux_50_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL not_4619_nl : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_re_mux_59_nl : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL not_4620_nl : STD_LOGIC;
  SIGNAL output_and_35_nl : STD_LOGIC;
  SIGNAL output_and_39_nl : STD_LOGIC;
  SIGNAL output_and_43_nl : STD_LOGIC;
  SIGNAL output_and_47_nl : STD_LOGIC;
  SIGNAL output_and_51_nl : STD_LOGIC;
  SIGNAL output_and_55_nl : STD_LOGIC;
  SIGNAL output_and_59_nl : STD_LOGIC;
  SIGNAL output_and_63_nl : STD_LOGIC;
  SIGNAL output_and_61_nl : STD_LOGIC;
  SIGNAL output_and_57_nl : STD_LOGIC;
  SIGNAL output_and_53_nl : STD_LOGIC;
  SIGNAL output_and_49_nl : STD_LOGIC;
  SIGNAL output_and_45_nl : STD_LOGIC;
  SIGNAL output_and_41_nl : STD_LOGIC;
  SIGNAL output_and_37_nl : STD_LOGIC;
  SIGNAL output_and_33_nl : STD_LOGIC;
  SIGNAL or_1659_nl : STD_LOGIC;
  SIGNAL nand_298_nl : STD_LOGIC;
  SIGNAL or_1661_nl : STD_LOGIC;
  SIGNAL nand_299_nl : STD_LOGIC;
  SIGNAL or_1663_nl : STD_LOGIC;
  SIGNAL nand_300_nl : STD_LOGIC;
  SIGNAL or_1665_nl : STD_LOGIC;
  SIGNAL nand_301_nl : STD_LOGIC;
  SIGNAL or_1669_nl : STD_LOGIC;
  SIGNAL or_1671_nl : STD_LOGIC;
  SIGNAL compute_sqrt_1_for_acc_1_nl : STD_LOGIC_VECTOR (40 DOWNTO 0);
  SIGNAL or_1860_nl : STD_LOGIC;
  SIGNAL compute_sqrt_for_acc_1_nl : STD_LOGIC_VECTOR (40 DOWNTO 0);
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_and_1_nl : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_2_acc_4_nl : STD_LOGIC_VECTOR (40 DOWNTO 0);
  SIGNAL QUANTIZE_ACTIVATION_LOOP_2_attention_abs_2_nand_nl : STD_LOGIC;
  SIGNAL attention_abs_2_mux_3_nl : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_nl : STD_LOGIC_VECTOR
      (25 DOWNTO 0);
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux_32_nl : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_3_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_1_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_4_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_2_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_5_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_3_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_6_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_4_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_7_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_5_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_8_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_6_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_9_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_7_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_17_nl : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_5_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_1_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_6_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_2_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_7_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_3_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_8_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_4_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_9_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_5_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_10_nl
      : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_6_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_11_nl
      : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_7_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_17_nl : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_mux_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_3_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_mux_1_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_4_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_mux_2_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_5_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_mux_3_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_6_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_mux_4_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_7_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_mux_5_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_8_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_mux_6_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_9_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_mux_7_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_1_nl
      : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_7_nl
      : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_25_nl
      : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_nl
      : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_6_nl
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_26_nl
      : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_27_nl
      : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_28_nl
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_16_nl
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_17_nl
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_18_nl
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_19_nl
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_20_nl
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_21_nl
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_22_nl
      : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_23_nl
      : STD_LOGIC;
  SIGNAL nand_378_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_nl : STD_LOGIC_VECTOR (55 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_nl : STD_LOGIC_VECTOR (55 DOWNTO 0);
  SIGNAL or_3014_nl : STD_LOGIC;
  SIGNAL or_3017_nl : STD_LOGIC;
  SIGNAL or_3019_nl : STD_LOGIC;
  SIGNAL or_3021_nl : STD_LOGIC;
  SIGNAL or_3022_nl : STD_LOGIC;
  SIGNAL or_3023_nl : STD_LOGIC;
  SIGNAL or_3024_nl : STD_LOGIC;
  SIGNAL or_3025_nl : STD_LOGIC;
  SIGNAL or_3027_nl : STD_LOGIC;
  SIGNAL or_3028_nl : STD_LOGIC;
  SIGNAL or_3029_nl : STD_LOGIC;
  SIGNAL or_3030_nl : STD_LOGIC;
  SIGNAL SF_LOOP_3_and_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_acc_nl : STD_LOGIC_VECTOR (23 DOWNTO
      0);
  SIGNAL QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_nl : STD_LOGIC_VECTOR (40 DOWNTO 0);
  SIGNAL QUANTIZE_ACTIVATION_LOOP_2_1_attention_abs_6_nand_nl : STD_LOGIC;
  SIGNAL attention_abs_6_mux_3_nl : STD_LOGIC_VECTOR (38 DOWNTO 0);
  SIGNAL QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_nl : STD_LOGIC_VECTOR
      (25 DOWNTO 0);
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_mux_32_nl : STD_LOGIC_VECTOR
      (23 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_3_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_1_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_4_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_2_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_5_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_3_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_6_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_4_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_7_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_5_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_8_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_6_nl : STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_9_nl :
      STD_LOGIC;
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_7_nl : STD_LOGIC;
  SIGNAL CACHE_UPDATE_LOOP_2_1_acc_2_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL attention_max_attn_fixed_t_1_acc_1_nl : STD_LOGIC_VECTOR (40 DOWNTO 0);
  SIGNAL CACHE_UPDATE_LOOP_2_acc_2_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL SOFTMAX_LOOP_3_acc_3_nl : STD_LOGIC_VECTOR (40 DOWNTO 0);
  SIGNAL mux_819_nl : STD_LOGIC;
  SIGNAL mux_817_nl : STD_LOGIC;
  SIGNAL mux_831_nl : STD_LOGIC;
  SIGNAL mux_830_nl : STD_LOGIC;
  SIGNAL mux_829_nl : STD_LOGIC;
  SIGNAL mux_828_nl : STD_LOGIC;
  SIGNAL mux_827_nl : STD_LOGIC;
  SIGNAL nand_257_nl : STD_LOGIC;
  SIGNAL or_1090_nl : STD_LOGIC;
  SIGNAL mux_826_nl : STD_LOGIC;
  SIGNAL mux_823_nl : STD_LOGIC;
  SIGNAL mux_822_nl : STD_LOGIC;
  SIGNAL mux_835_nl : STD_LOGIC;
  SIGNAL mux_833_nl : STD_LOGIC;
  SIGNAL mux_837_nl : STD_LOGIC;
  SIGNAL and_1498_nl : STD_LOGIC;
  SIGNAL nor_897_nl : STD_LOGIC;
  SIGNAL and_337_nl : STD_LOGIC;
  SIGNAL mux_858_nl : STD_LOGIC;
  SIGNAL mux_867_nl : STD_LOGIC;
  SIGNAL nand_262_nl : STD_LOGIC;
  SIGNAL mux_866_nl : STD_LOGIC;
  SIGNAL and_344_nl : STD_LOGIC;
  SIGNAL or_3142_nl : STD_LOGIC;
  SIGNAL mux_865_nl : STD_LOGIC;
  SIGNAL or_1827_nl : STD_LOGIC;
  SIGNAL mux_904_nl : STD_LOGIC;
  SIGNAL nand_44_nl : STD_LOGIC;
  SIGNAL mux_903_nl : STD_LOGIC;
  SIGNAL mux_953_nl : STD_LOGIC;
  SIGNAL or_3149_nl : STD_LOGIC;
  SIGNAL or_3150_nl : STD_LOGIC;
  SIGNAL nor_923_nl : STD_LOGIC;
  SIGNAL nand_264_nl : STD_LOGIC;
  SIGNAL or_1910_nl : STD_LOGIC;
  SIGNAL or_1912_nl : STD_LOGIC;
  SIGNAL or_3073_nl : STD_LOGIC;
  SIGNAL mux_1026_nl : STD_LOGIC;
  SIGNAL mux_1028_nl : STD_LOGIC;
  SIGNAL or_1976_nl : STD_LOGIC;
  SIGNAL or_1974_nl : STD_LOGIC;
  SIGNAL mux_1149_nl : STD_LOGIC;
  SIGNAL mux_1148_nl : STD_LOGIC;
  SIGNAL mux_1162_nl : STD_LOGIC;
  SIGNAL mux_1161_nl : STD_LOGIC;
  SIGNAL mux_1160_nl : STD_LOGIC;
  SIGNAL mux_1159_nl : STD_LOGIC;
  SIGNAL mux_1158_nl : STD_LOGIC;
  SIGNAL mux_1157_nl : STD_LOGIC;
  SIGNAL mux_1156_nl : STD_LOGIC;
  SIGNAL mux_1155_nl : STD_LOGIC;
  SIGNAL mux_1154_nl : STD_LOGIC;
  SIGNAL mux_1153_nl : STD_LOGIC;
  SIGNAL mux_1152_nl : STD_LOGIC;
  SIGNAL mux_1249_nl : STD_LOGIC;
  SIGNAL mux_1311_nl : STD_LOGIC;
  SIGNAL or_2235_nl : STD_LOGIC;
  SIGNAL mux_1313_nl : STD_LOGIC;
  SIGNAL nor_930_nl : STD_LOGIC;
  SIGNAL mux_1312_nl : STD_LOGIC;
  SIGNAL and_443_nl : STD_LOGIC;
  SIGNAL mux_1400_nl : STD_LOGIC;
  SIGNAL mux_1399_nl : STD_LOGIC;
  SIGNAL mux_1398_nl : STD_LOGIC;
  SIGNAL mux_1396_nl : STD_LOGIC;
  SIGNAL and_1616_nl : STD_LOGIC;
  SIGNAL mux_1395_nl : STD_LOGIC;
  SIGNAL mux_1394_nl : STD_LOGIC;
  SIGNAL or_2296_nl : STD_LOGIC;
  SIGNAL mux_1406_nl : STD_LOGIC;
  SIGNAL or_2309_nl : STD_LOGIC;
  SIGNAL mux_1405_nl : STD_LOGIC;
  SIGNAL mux_1404_nl : STD_LOGIC;
  SIGNAL or_1049_nl : STD_LOGIC;
  SIGNAL or_2322_nl : STD_LOGIC;
  SIGNAL mux_1422_nl : STD_LOGIC;
  SIGNAL and_1303_nl : STD_LOGIC;
  SIGNAL mux_1425_nl : STD_LOGIC;
  SIGNAL mux_1424_nl : STD_LOGIC;
  SIGNAL mux_1423_nl : STD_LOGIC;
  SIGNAL mux_1427_nl : STD_LOGIC;
  SIGNAL or_2328_nl : STD_LOGIC;
  SIGNAL mux_1436_nl : STD_LOGIC;
  SIGNAL nor_938_nl : STD_LOGIC;
  SIGNAL mux_1435_nl : STD_LOGIC;
  SIGNAL nor_939_nl : STD_LOGIC;
  SIGNAL mux_1450_nl : STD_LOGIC;
  SIGNAL mux_1449_nl : STD_LOGIC;
  SIGNAL mux_137_nl : STD_LOGIC;
  SIGNAL mux_1942_nl : STD_LOGIC;
  SIGNAL nor_946_nl : STD_LOGIC;
  SIGNAL mux_1944_nl : STD_LOGIC;
  SIGNAL or_2744_nl : STD_LOGIC;
  SIGNAL mux_2035_nl : STD_LOGIC;
  SIGNAL or_2746_nl : STD_LOGIC;
  SIGNAL mux_2066_nl : STD_LOGIC;
  SIGNAL mux_2085_nl : STD_LOGIC;
  SIGNAL or_2784_nl : STD_LOGIC;
  SIGNAL mux_2113_nl : STD_LOGIC;
  SIGNAL mux_2112_nl : STD_LOGIC;
  SIGNAL mux_2111_nl : STD_LOGIC;
  SIGNAL nor_953_nl : STD_LOGIC;
  SIGNAL nor_954_nl : STD_LOGIC;
  SIGNAL nor_955_nl : STD_LOGIC;
  SIGNAL mux_2110_nl : STD_LOGIC;
  SIGNAL or_2833_nl : STD_LOGIC;
  SIGNAL nor_956_nl : STD_LOGIC;
  SIGNAL mux_2115_nl : STD_LOGIC;
  SIGNAL mux_2117_nl : STD_LOGIC;
  SIGNAL nor_957_nl : STD_LOGIC;
  SIGNAL mux_2118_nl : STD_LOGIC;
  SIGNAL mux_2152_nl : STD_LOGIC;
  SIGNAL mux_2151_nl : STD_LOGIC;
  SIGNAL mux_2150_nl : STD_LOGIC;
  SIGNAL mux_2149_nl : STD_LOGIC;
  SIGNAL mux_2148_nl : STD_LOGIC;
  SIGNAL mux_2147_nl : STD_LOGIC;
  SIGNAL nand_286_nl : STD_LOGIC;
  SIGNAL or_2872_nl : STD_LOGIC;
  SIGNAL mux_2145_nl : STD_LOGIC;
  SIGNAL nand_101_nl : STD_LOGIC;
  SIGNAL or_2869_nl : STD_LOGIC;
  SIGNAL mux_2144_nl : STD_LOGIC;
  SIGNAL or_2868_nl : STD_LOGIC;
  SIGNAL mux_2143_nl : STD_LOGIC;
  SIGNAL mux_2142_nl : STD_LOGIC;
  SIGNAL or_2866_nl : STD_LOGIC;
  SIGNAL mux_2175_nl : STD_LOGIC;
  SIGNAL mux_2174_nl : STD_LOGIC;
  SIGNAL mux_2173_nl : STD_LOGIC;
  SIGNAL mux_2172_nl : STD_LOGIC;
  SIGNAL mux_2171_nl : STD_LOGIC;
  SIGNAL mux_2170_nl : STD_LOGIC;
  SIGNAL or_2901_nl : STD_LOGIC;
  SIGNAL mux_2169_nl : STD_LOGIC;
  SIGNAL mux_2168_nl : STD_LOGIC;
  SIGNAL and_1544_nl : STD_LOGIC;
  SIGNAL mux_2165_nl : STD_LOGIC;
  SIGNAL mux_2164_nl : STD_LOGIC;
  SIGNAL mux_2162_nl : STD_LOGIC;
  SIGNAL mux_2161_nl : STD_LOGIC;
  SIGNAL mux_2160_nl : STD_LOGIC;
  SIGNAL or_2897_nl : STD_LOGIC;
  SIGNAL or_2894_nl : STD_LOGIC;
  SIGNAL or_2890_nl : STD_LOGIC;
  SIGNAL mux_2251_nl : STD_LOGIC;
  SIGNAL and_1546_nl : STD_LOGIC;
  SIGNAL nor_968_nl : STD_LOGIC;
  SIGNAL or_3055_nl : STD_LOGIC;
  SIGNAL or_3058_nl : STD_LOGIC;
  SIGNAL mux_2255_nl : STD_LOGIC;
  SIGNAL mux_2254_nl : STD_LOGIC;
  SIGNAL mux_2253_nl : STD_LOGIC;
  SIGNAL or_1418_nl : STD_LOGIC;
  SIGNAL nand_295_nl : STD_LOGIC;
  SIGNAL mux_2259_nl : STD_LOGIC;
  SIGNAL and_1550_nl : STD_LOGIC;
  SIGNAL nor_969_nl : STD_LOGIC;
  SIGNAL mux_869_nl : STD_LOGIC;
  SIGNAL mux_868_nl : STD_LOGIC;
  SIGNAL mux_1010_nl : STD_LOGIC;
  SIGNAL mux_1009_nl : STD_LOGIC;
  SIGNAL mux_1008_nl : STD_LOGIC;
  SIGNAL mux_1007_nl : STD_LOGIC;
  SIGNAL nor_999_nl : STD_LOGIC;
  SIGNAL mux_1006_nl : STD_LOGIC;
  SIGNAL mux_1005_nl : STD_LOGIC;
  SIGNAL nand_322_nl : STD_LOGIC;
  SIGNAL nor_1001_nl : STD_LOGIC;
  SIGNAL mux_1004_nl : STD_LOGIC;
  SIGNAL mux_1003_nl : STD_LOGIC;
  SIGNAL or_1952_nl : STD_LOGIC;
  SIGNAL or_1950_nl : STD_LOGIC;
  SIGNAL mux_1002_nl : STD_LOGIC;
  SIGNAL mux_1001_nl : STD_LOGIC;
  SIGNAL nand_323_nl : STD_LOGIC;
  SIGNAL mux_999_nl : STD_LOGIC;
  SIGNAL mux_998_nl : STD_LOGIC;
  SIGNAL nand_325_nl : STD_LOGIC;
  SIGNAL mux_997_nl : STD_LOGIC;
  SIGNAL or_1944_nl : STD_LOGIC;
  SIGNAL mux_996_nl : STD_LOGIC;
  SIGNAL mux_995_nl : STD_LOGIC;
  SIGNAL mux_994_nl : STD_LOGIC;
  SIGNAL mux_993_nl : STD_LOGIC;
  SIGNAL or_1943_nl : STD_LOGIC;
  SIGNAL mux_992_nl : STD_LOGIC;
  SIGNAL mux_991_nl : STD_LOGIC;
  SIGNAL or_1940_nl : STD_LOGIC;
  SIGNAL mux_990_nl : STD_LOGIC;
  SIGNAL mux_989_nl : STD_LOGIC;
  SIGNAL mux_988_nl : STD_LOGIC;
  SIGNAL mux_987_nl : STD_LOGIC;
  SIGNAL or_1939_nl : STD_LOGIC;
  SIGNAL or_1938_nl : STD_LOGIC;
  SIGNAL or_1937_nl : STD_LOGIC;
  SIGNAL or_1934_nl : STD_LOGIC;
  SIGNAL or_1933_nl : STD_LOGIC;
  SIGNAL mux_986_nl : STD_LOGIC;
  SIGNAL or_1932_nl : STD_LOGIC;
  SIGNAL or_1931_nl : STD_LOGIC;
  SIGNAL mux_1025_nl : STD_LOGIC;
  SIGNAL mux_1024_nl : STD_LOGIC;
  SIGNAL nor_1019_nl : STD_LOGIC;
  SIGNAL mux_1023_nl : STD_LOGIC;
  SIGNAL mux_1022_nl : STD_LOGIC;
  SIGNAL mux_1021_nl : STD_LOGIC;
  SIGNAL nor_1020_nl : STD_LOGIC;
  SIGNAL nor_1021_nl : STD_LOGIC;
  SIGNAL mux_1020_nl : STD_LOGIC;
  SIGNAL nor_1022_nl : STD_LOGIC;
  SIGNAL mux_1019_nl : STD_LOGIC;
  SIGNAL nor_1023_nl : STD_LOGIC;
  SIGNAL nor_1024_nl : STD_LOGIC;
  SIGNAL mux_1032_nl : STD_LOGIC;
  SIGNAL nand_49_nl : STD_LOGIC;
  SIGNAL mux_1031_nl : STD_LOGIC;
  SIGNAL mux_1030_nl : STD_LOGIC;
  SIGNAL mux_1029_nl : STD_LOGIC;
  SIGNAL mux_1078_nl : STD_LOGIC;
  SIGNAL nor_1031_nl : STD_LOGIC;
  SIGNAL nand_330_nl : STD_LOGIC;
  SIGNAL mux_1076_nl : STD_LOGIC;
  SIGNAL nor_1032_nl : STD_LOGIC;
  SIGNAL nor_1033_nl : STD_LOGIC;
  SIGNAL mux_1073_nl : STD_LOGIC;
  SIGNAL or_2022_nl : STD_LOGIC;
  SIGNAL mux_1077_nl : STD_LOGIC;
  SIGNAL mux_1075_nl : STD_LOGIC;
  SIGNAL or_2019_nl : STD_LOGIC;
  SIGNAL mux_1088_nl : STD_LOGIC;
  SIGNAL nand_52_nl : STD_LOGIC;
  SIGNAL mux_1086_nl : STD_LOGIC;
  SIGNAL mux_1085_nl : STD_LOGIC;
  SIGNAL or_2038_nl : STD_LOGIC;
  SIGNAL mux_1083_nl : STD_LOGIC;
  SIGNAL mux_1082_nl : STD_LOGIC;
  SIGNAL nand_332_nl : STD_LOGIC;
  SIGNAL nand_51_nl : STD_LOGIC;
  SIGNAL mux_1081_nl : STD_LOGIC;
  SIGNAL nor_1035_nl : STD_LOGIC;
  SIGNAL nor_1036_nl : STD_LOGIC;
  SIGNAL or_2034_nl : STD_LOGIC;
  SIGNAL mux_1080_nl : STD_LOGIC;
  SIGNAL mux_1091_nl : STD_LOGIC;
  SIGNAL or_2041_nl : STD_LOGIC;
  SIGNAL mux_1090_nl : STD_LOGIC;
  SIGNAL or_2039_nl : STD_LOGIC;
  SIGNAL mux_1111_nl : STD_LOGIC;
  SIGNAL or_2070_nl : STD_LOGIC;
  SIGNAL mux_1110_nl : STD_LOGIC;
  SIGNAL or_2068_nl : STD_LOGIC;
  SIGNAL mux_1131_nl : STD_LOGIC;
  SIGNAL mux_1130_nl : STD_LOGIC;
  SIGNAL mux_1129_nl : STD_LOGIC;
  SIGNAL mux_1128_nl : STD_LOGIC;
  SIGNAL mux_1127_nl : STD_LOGIC;
  SIGNAL mux_1126_nl : STD_LOGIC;
  SIGNAL mux_1123_nl : STD_LOGIC;
  SIGNAL mux_1121_nl : STD_LOGIC;
  SIGNAL or_2095_nl : STD_LOGIC;
  SIGNAL or_2110_nl : STD_LOGIC;
  SIGNAL mux_1196_nl : STD_LOGIC;
  SIGNAL mux_1195_nl : STD_LOGIC;
  SIGNAL mux_1194_nl : STD_LOGIC;
  SIGNAL mux_1193_nl : STD_LOGIC;
  SIGNAL mux_1192_nl : STD_LOGIC;
  SIGNAL mux_1191_nl : STD_LOGIC;
  SIGNAL mux_1190_nl : STD_LOGIC;
  SIGNAL mux_1189_nl : STD_LOGIC;
  SIGNAL mux_1188_nl : STD_LOGIC;
  SIGNAL mux_1186_nl : STD_LOGIC;
  SIGNAL mux_1184_nl : STD_LOGIC;
  SIGNAL mux_1182_nl : STD_LOGIC;
  SIGNAL mux_1181_nl : STD_LOGIC;
  SIGNAL mux_1180_nl : STD_LOGIC;
  SIGNAL or_2121_nl : STD_LOGIC;
  SIGNAL and_1593_nl : STD_LOGIC;
  SIGNAL or_2132_nl : STD_LOGIC;
  SIGNAL mux_1206_nl : STD_LOGIC;
  SIGNAL mux_1205_nl : STD_LOGIC;
  SIGNAL nor_1043_nl : STD_LOGIC;
  SIGNAL and_1595_nl : STD_LOGIC;
  SIGNAL mux_1204_nl : STD_LOGIC;
  SIGNAL mux_1203_nl : STD_LOGIC;
  SIGNAL or_2130_nl : STD_LOGIC;
  SIGNAL mux_1202_nl : STD_LOGIC;
  SIGNAL or_3166_nl : STD_LOGIC;
  SIGNAL mux_1201_nl : STD_LOGIC;
  SIGNAL or_2129_nl : STD_LOGIC;
  SIGNAL mux_1200_nl : STD_LOGIC;
  SIGNAL mux_1199_nl : STD_LOGIC;
  SIGNAL or_2127_nl : STD_LOGIC;
  SIGNAL mux_1198_nl : STD_LOGIC;
  SIGNAL or_2126_nl : STD_LOGIC;
  SIGNAL nor_1325_nl : STD_LOGIC;
  SIGNAL mux_1273_nl : STD_LOGIC;
  SIGNAL mux_1272_nl : STD_LOGIC;
  SIGNAL mux_1271_nl : STD_LOGIC;
  SIGNAL mux_1270_nl : STD_LOGIC;
  SIGNAL or_2184_nl : STD_LOGIC;
  SIGNAL nor_1050_nl : STD_LOGIC;
  SIGNAL mux_1269_nl : STD_LOGIC;
  SIGNAL mux_1268_nl : STD_LOGIC;
  SIGNAL mux_1267_nl : STD_LOGIC;
  SIGNAL mux_1266_nl : STD_LOGIC;
  SIGNAL mux_1265_nl : STD_LOGIC;
  SIGNAL nor_1326_nl : STD_LOGIC;
  SIGNAL nor_1327_nl : STD_LOGIC;
  SIGNAL mux_1264_nl : STD_LOGIC;
  SIGNAL mux_1263_nl : STD_LOGIC;
  SIGNAL nor_1328_nl : STD_LOGIC;
  SIGNAL nor_1329_nl : STD_LOGIC;
  SIGNAL mux_1262_nl : STD_LOGIC;
  SIGNAL nor_1330_nl : STD_LOGIC;
  SIGNAL nor_1331_nl : STD_LOGIC;
  SIGNAL mux_1276_nl : STD_LOGIC;
  SIGNAL mux_1275_nl : STD_LOGIC;
  SIGNAL nor_1054_nl : STD_LOGIC;
  SIGNAL nor_1055_nl : STD_LOGIC;
  SIGNAL mux_1280_nl : STD_LOGIC;
  SIGNAL or_3169_nl : STD_LOGIC;
  SIGNAL mux_1279_nl : STD_LOGIC;
  SIGNAL or_2199_nl : STD_LOGIC;
  SIGNAL or_2198_nl : STD_LOGIC;
  SIGNAL or_3170_nl : STD_LOGIC;
  SIGNAL mux_1278_nl : STD_LOGIC;
  SIGNAL or_2195_nl : STD_LOGIC;
  SIGNAL mux_1277_nl : STD_LOGIC;
  SIGNAL or_2193_nl : STD_LOGIC;
  SIGNAL mux_1284_nl : STD_LOGIC;
  SIGNAL mux_1283_nl : STD_LOGIC;
  SIGNAL and_601_nl : STD_LOGIC;
  SIGNAL nor_1060_nl : STD_LOGIC;
  SIGNAL mux_1282_nl : STD_LOGIC;
  SIGNAL or_2203_nl : STD_LOGIC;
  SIGNAL nor_1102_nl : STD_LOGIC;
  SIGNAL and_1635_nl : STD_LOGIC;
  SIGNAL mux_1402_nl : STD_LOGIC;
  SIGNAL mux_1401_nl : STD_LOGIC;
  SIGNAL nor_1099_nl : STD_LOGIC;
  SIGNAL nor_1100_nl : STD_LOGIC;
  SIGNAL nor_1101_nl : STD_LOGIC;
  SIGNAL mux_1409_nl : STD_LOGIC;
  SIGNAL mux_1408_nl : STD_LOGIC;
  SIGNAL mux_1407_nl : STD_LOGIC;
  SIGNAL mux_1448_nl : STD_LOGIC;
  SIGNAL and_1642_nl : STD_LOGIC;
  SIGNAL mux_1447_nl : STD_LOGIC;
  SIGNAL nor_1111_nl : STD_LOGIC;
  SIGNAL mux_1446_nl : STD_LOGIC;
  SIGNAL mux_1445_nl : STD_LOGIC;
  SIGNAL mux_1444_nl : STD_LOGIC;
  SIGNAL mux_1443_nl : STD_LOGIC;
  SIGNAL mux_1442_nl : STD_LOGIC;
  SIGNAL and_1644_nl : STD_LOGIC;
  SIGNAL mux_1464_nl : STD_LOGIC;
  SIGNAL nor_1118_nl : STD_LOGIC;
  SIGNAL nor_1119_nl : STD_LOGIC;
  SIGNAL mux_1463_nl : STD_LOGIC;
  SIGNAL nor_1120_nl : STD_LOGIC;
  SIGNAL mux_1462_nl : STD_LOGIC;
  SIGNAL nor_1121_nl : STD_LOGIC;
  SIGNAL mux_1461_nl : STD_LOGIC;
  SIGNAL or_2363_nl : STD_LOGIC;
  SIGNAL or_2362_nl : STD_LOGIC;
  SIGNAL mux_1460_nl : STD_LOGIC;
  SIGNAL mux_1459_nl : STD_LOGIC;
  SIGNAL nor_1122_nl : STD_LOGIC;
  SIGNAL nor_1123_nl : STD_LOGIC;
  SIGNAL mux_1458_nl : STD_LOGIC;
  SIGNAL nor_1124_nl : STD_LOGIC;
  SIGNAL nor_1125_nl : STD_LOGIC;
  SIGNAL mux_1474_nl : STD_LOGIC;
  SIGNAL mux_1473_nl : STD_LOGIC;
  SIGNAL nor_1129_nl : STD_LOGIC;
  SIGNAL nor_1130_nl : STD_LOGIC;
  SIGNAL and_1646_nl : STD_LOGIC;
  SIGNAL mux_1472_nl : STD_LOGIC;
  SIGNAL nor_1126_nl : STD_LOGIC;
  SIGNAL mux_1471_nl : STD_LOGIC;
  SIGNAL nor_1127_nl : STD_LOGIC;
  SIGNAL nor_1128_nl : STD_LOGIC;
  SIGNAL mux_1470_nl : STD_LOGIC;
  SIGNAL mux_1469_nl : STD_LOGIC;
  SIGNAL nor_1131_nl : STD_LOGIC;
  SIGNAL nor_1132_nl : STD_LOGIC;
  SIGNAL mux_1468_nl : STD_LOGIC;
  SIGNAL mux_1467_nl : STD_LOGIC;
  SIGNAL nor_1133_nl : STD_LOGIC;
  SIGNAL nor_1134_nl : STD_LOGIC;
  SIGNAL nor_1135_nl : STD_LOGIC;
  SIGNAL mux_1586_nl : STD_LOGIC;
  SIGNAL or_2499_nl : STD_LOGIC;
  SIGNAL mux_1592_nl : STD_LOGIC;
  SIGNAL nand_359_nl : STD_LOGIC;
  SIGNAL mux_1594_nl : STD_LOGIC;
  SIGNAL mux_2262_nl : STD_LOGIC;
  SIGNAL mux_1595_nl : STD_LOGIC;
  SIGNAL mux_1593_nl : STD_LOGIC;
  SIGNAL mux_1596_nl : STD_LOGIC;
  SIGNAL mux_1598_nl : STD_LOGIC;
  SIGNAL mux_1597_nl : STD_LOGIC;
  SIGNAL and_1659_nl : STD_LOGIC;
  SIGNAL mux_1599_nl : STD_LOGIC;
  SIGNAL mux_1607_nl : STD_LOGIC;
  SIGNAL mux_1606_nl : STD_LOGIC;
  SIGNAL nor_1160_nl : STD_LOGIC;
  SIGNAL mux_1605_nl : STD_LOGIC;
  SIGNAL nand_361_nl : STD_LOGIC;
  SIGNAL nand_362_nl : STD_LOGIC;
  SIGNAL mux_1604_nl : STD_LOGIC;
  SIGNAL nor_1161_nl : STD_LOGIC;
  SIGNAL mux_1603_nl : STD_LOGIC;
  SIGNAL nor_1162_nl : STD_LOGIC;
  SIGNAL nor_1163_nl : STD_LOGIC;
  SIGNAL mux_1602_nl : STD_LOGIC;
  SIGNAL nor_1164_nl : STD_LOGIC;
  SIGNAL nor_1165_nl : STD_LOGIC;
  SIGNAL mux_1601_nl : STD_LOGIC;
  SIGNAL mux_1608_nl : STD_LOGIC;
  SIGNAL and_1667_nl : STD_LOGIC;
  SIGNAL mux_1610_nl : STD_LOGIC;
  SIGNAL and_1666_nl : STD_LOGIC;
  SIGNAL nor_1169_nl : STD_LOGIC;
  SIGNAL and_1668_nl : STD_LOGIC;
  SIGNAL mux_1609_nl : STD_LOGIC;
  SIGNAL nor_1170_nl : STD_LOGIC;
  SIGNAL nor_1171_nl : STD_LOGIC;
  SIGNAL mux_1615_nl : STD_LOGIC;
  SIGNAL mux_1614_nl : STD_LOGIC;
  SIGNAL or_2541_nl : STD_LOGIC;
  SIGNAL or_3189_nl : STD_LOGIC;
  SIGNAL mux_2060_nl : STD_LOGIC;
  SIGNAL or_2762_nl : STD_LOGIC;
  SIGNAL mux_2069_nl : STD_LOGIC;
  SIGNAL or_2768_nl : STD_LOGIC;
  SIGNAL mux_2138_nl : STD_LOGIC;
  SIGNAL and_1778_nl : STD_LOGIC;
  SIGNAL mux_2137_nl : STD_LOGIC;
  SIGNAL mux_2136_nl : STD_LOGIC;
  SIGNAL or_1238_nl : STD_LOGIC;
  SIGNAL nor_1234_nl : STD_LOGIC;
  SIGNAL mux_2140_nl : STD_LOGIC;
  SIGNAL mux_2135_nl : STD_LOGIC;
  SIGNAL mux_2134_nl : STD_LOGIC;
  SIGNAL mux_2133_nl : STD_LOGIC;
  SIGNAL mux_2132_nl : STD_LOGIC;
  SIGNAL and_1780_nl : STD_LOGIC;
  SIGNAL nor_1261_nl : STD_LOGIC;
  SIGNAL mux_2191_nl : STD_LOGIC;
  SIGNAL mux_2186_nl : STD_LOGIC;
  SIGNAL mux_2185_nl : STD_LOGIC;
  SIGNAL mux_2184_nl : STD_LOGIC;
  SIGNAL mux_2183_nl : STD_LOGIC;
  SIGNAL nor_1299_nl : STD_LOGIC;
  SIGNAL mux_2219_nl : STD_LOGIC;
  SIGNAL mux_2214_nl : STD_LOGIC;
  SIGNAL mux_2213_nl : STD_LOGIC;
  SIGNAL mux_2212_nl : STD_LOGIC;
  SIGNAL mux_2211_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_l_mux1h_6_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_4_l_mux1h_8_nl : STD_LOGIC;
  SIGNAL QUANTIZE_ACTIVATION_LOOP_1_1_max_val_asn_GEMM_3D_FLOAT_LOOP_4_l_2_operator_40_24_true_AC_TRN_AC_WRAP_or_nl
      : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_mux1h_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_or_nl : STD_LOGIC;
  SIGNAL compute_sqrt_for_acc_3_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_2_and_35_nl : STD_LOGIC;
  SIGNAL nor_658_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_and_35_nl : STD_LOGIC;
  SIGNAL mux_1260_nl : STD_LOGIC;
  SIGNAL mux_1259_nl : STD_LOGIC;
  SIGNAL mux_1258_nl : STD_LOGIC;
  SIGNAL mux_1257_nl : STD_LOGIC;
  SIGNAL mux_1256_nl : STD_LOGIC;
  SIGNAL mux_1255_nl : STD_LOGIC;
  SIGNAL mux_1254_nl : STD_LOGIC;
  SIGNAL mux_1253_nl : STD_LOGIC;
  SIGNAL mux_1252_nl : STD_LOGIC;
  SIGNAL or_2167_nl : STD_LOGIC;
  SIGNAL mux_1251_nl : STD_LOGIC;
  SIGNAL mux_1247_nl : STD_LOGIC;
  SIGNAL mux_1246_nl : STD_LOGIC;
  SIGNAL mux_1244_nl : STD_LOGIC;
  SIGNAL mux_1243_nl : STD_LOGIC;
  SIGNAL or_3075_nl : STD_LOGIC;
  SIGNAL mux_1242_nl : STD_LOGIC;
  SIGNAL mux_1241_nl : STD_LOGIC;
  SIGNAL nor_374_nl : STD_LOGIC;
  SIGNAL mux_1239_nl : STD_LOGIC;
  SIGNAL or_2162_nl : STD_LOGIC;
  SIGNAL mux_1261_nl : STD_LOGIC;
  SIGNAL nor_1048_nl : STD_LOGIC;
  SIGNAL and_1603_nl : STD_LOGIC;
  SIGNAL and_1256_nl : STD_LOGIC;
  SIGNAL and_1257_nl : STD_LOGIC;
  SIGNAL mux_2247_nl : STD_LOGIC;
  SIGNAL mux_2246_nl : STD_LOGIC;
  SIGNAL nor_1318_nl : STD_LOGIC;
  SIGNAL CACHE_UPDATE_LOOP_3_mux_3_nl : STD_LOGIC_VECTOR (39 DOWNTO 0);
  SIGNAL and_369_nl : STD_LOGIC;
  SIGNAL TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL CACHE_UPDATE_LOOP_3_acc_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL CACHE_UPDATE_LOOP_3_1_CACHE_UPDATE_LOOP_3_1_mux_nl : STD_LOGIC_VECTOR (23
      DOWNTO 0);
  SIGNAL CACHE_UPDATE_LOOP_3_1_mux_2_nl : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL CACHE_UPDATE_LOOP_3_1_CACHE_UPDATE_LOOP_3_1_mux_1_nl : STD_LOGIC_VECTOR
      (15 DOWNTO 0);
  SIGNAL CACHE_UPDATE_LOOP_3_1_mux_3_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_4_1_acc_13_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL GEMM_3D_FLOAT_LOOP_4_acc_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL mux_2299_nl : STD_LOGIC;
  SIGNAL nor_1345_nl : STD_LOGIC;
  SIGNAL nor_1346_nl : STD_LOGIC;
  SIGNAL mux_2288_nl : STD_LOGIC;
  SIGNAL nor_1378_nl : STD_LOGIC;
  SIGNAL nor_1379_nl : STD_LOGIC;
  SIGNAL mux_2292_nl : STD_LOGIC;
  SIGNAL or_3261_nl : STD_LOGIC;
  SIGNAL mux_2291_nl : STD_LOGIC;
  SIGNAL mux_2290_nl : STD_LOGIC;
  SIGNAL or_3235_nl : STD_LOGIC;
  SIGNAL mux_2267_nl : STD_LOGIC;
  SIGNAL mux_2266_nl : STD_LOGIC;
  SIGNAL nor_1348_nl : STD_LOGIC;
  SIGNAL mux_2268_nl : STD_LOGIC;
  SIGNAL nor_1350_nl : STD_LOGIC;
  SIGNAL mux_2270_nl : STD_LOGIC;
  SIGNAL nand_394_nl : STD_LOGIC;
  SIGNAL mux_2287_nl : STD_LOGIC;
  SIGNAL nor_1368_nl : STD_LOGIC;
  SIGNAL mux_2286_nl : STD_LOGIC;
  SIGNAL nand_398_nl : STD_LOGIC;
  SIGNAL nor_1369_nl : STD_LOGIC;
  SIGNAL CACHE_UPDATE_LOOP_3_mux1h_6_nl : STD_LOGIC;
  SIGNAL CACHE_UPDATE_LOOP_3_mux1h_7_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_1_GEMM_3D_FLOAT_LOOP_1_mux_2_nl : STD_LOGIC;
  SIGNAL GEMM_3D_FLOAT_LOOP_1_GEMM_3D_FLOAT_LOOP_1_mux_3_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_APPLY_ROTARY_POS_EMB_LOOP_6_or_8_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_36_nl : STD_LOGIC_VECTOR (12 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_37_nl : STD_LOGIC_VECTOR (23 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_38_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_39_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_40_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_41_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_42_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_43_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_44_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_45_nl : STD_LOGIC;
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_46_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_and_14_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_134_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_and_15_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_135_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_136_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_137_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_138_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_139_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_140_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_141_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_and_16_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_142_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_and_17_nl : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_143_nl : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_and_18_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_144_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL not_5114_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_3_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_145_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_4_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_146_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_and_19_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_147_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_5_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_148_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_149_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_and_20_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_150_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_or_13_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_151_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_152_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_or_14_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_153_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_1_1_mux1h_154_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_1_1_or_15_nl : STD_LOGIC;
  SIGNAL TRANSPOSE_LAST_TWO_DIMS_LOOP_3_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_mux_2_nl :
      STD_LOGIC;
  SIGNAL TRANSPOSE_LAST_TWO_DIMS_LOOP_3_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_mux_3_nl :
      STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_mux_1_nl : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL RMS_NORM_LOOP_2_2_or_1_nl : STD_LOGIC;
  SIGNAL mux_2300_nl : STD_LOGIC;
  SIGNAL mux_2301_nl : STD_LOGIC;
  SIGNAL mux_2302_nl : STD_LOGIC;
  SIGNAL nor_1397_nl : STD_LOGIC;
  SIGNAL mux_2303_nl : STD_LOGIC;
  SIGNAL nor_1398_nl : STD_LOGIC;
  SIGNAL and_2128_nl : STD_LOGIC;
  SIGNAL mul_3_nl : STD_LOGIC_VECTOR (71 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_2_2_mux_28_nl : STD_LOGIC_VECTOR (52 DOWNTO 0);
  SIGNAL and_2129_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_21_nl : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_22_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_23_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_22_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_23_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_24_nl : STD_LOGIC;
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_25_nl : STD_LOGIC;
  SIGNAL RMS_NORM_LOOP_2_2_mux_29_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL RMS_NORM_LOOP_2_2_mux_30_nl : STD_LOGIC;
  SIGNAL SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a : STD_LOGIC_VECTOR (55 DOWNTO
      0);
  SIGNAL SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z_1 : STD_LOGIC_VECTOR (55 DOWNTO
      0);

  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a
      : STD_LOGIC_VECTOR (71 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b
      : STD_LOGIC_VECTOR (59 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z_1
      : STD_LOGIC_VECTOR (71 DOWNTO 0);

  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_1 : STD_LOGIC_VECTOR (39
      DOWNTO 0);

  SIGNAL CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_rg_addr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_rg_data_out : STD_LOGIC_VECTOR
      (19 DOWNTO 0);

  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_rg_addr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_rg_data_out
      : STD_LOGIC_VECTOR (7 DOWNTO 0);

  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_rg_addr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_rg_data_out
      : STD_LOGIC_VECTOR (7 DOWNTO 0);

  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_rg_addr :
      STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_rg_data_out
      : STD_LOGIC_VECTOR (14 DOWNTO 0);

  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_rg_addr :
      STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_rg_data_out
      : STD_LOGIC_VECTOR (12 DOWNTO 0);

  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_rg_addr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_rg_data_out
      : STD_LOGIC_VECTOR (7 DOWNTO 0);

  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_rg_addr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_rg_data_out
      : STD_LOGIC_VECTOR (7 DOWNTO 0);

  SIGNAL CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_rg_addr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_rg_data_out : STD_LOGIC_VECTOR
      (18 DOWNTO 0);

  COMPONENT dut_core_strm_in_rsci
    PORT(
      strm_in_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      strm_in_rsc_vld : IN STD_LOGIC;
      strm_in_rsc_rdy : OUT STD_LOGIC;
      strm_in_rsci_oswt : IN STD_LOGIC;
      strm_in_rsci_wen_comp : OUT STD_LOGIC;
      strm_in_rsci_idat_mxwt : OUT STD_LOGIC_VECTOR (29 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL dut_core_strm_in_rsci_inst_strm_in_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL dut_core_strm_in_rsci_inst_strm_in_rsci_idat_mxwt : STD_LOGIC_VECTOR (29
      DOWNTO 0);

  COMPONENT dut_core_strm_out_rsci
    PORT(
      strm_out_rsc_dat : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      strm_out_rsc_vld : OUT STD_LOGIC;
      strm_out_rsc_rdy : IN STD_LOGIC;
      strm_out_rsci_oswt : IN STD_LOGIC;
      strm_out_rsci_wen_comp : OUT STD_LOGIC;
      strm_out_rsci_idat : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL dut_core_strm_out_rsci_inst_strm_out_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL dut_core_strm_out_rsci_inst_strm_out_rsci_idat : STD_LOGIC_VECTOR (31 DOWNTO
      0);

  COMPONENT dut_core_staller
    PORT(
      en : IN STD_LOGIC;
      core_wen1 : OUT STD_LOGIC;
      strm_in_rsci_wen_comp : IN STD_LOGIC;
      strm_out_rsci_wen_comp : IN STD_LOGIC;
      attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 : OUT STD_LOGIC
    );
  END COMPONENT;
  COMPONENT dut_core_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      rms_norm_16_div_cmp_z : IN STD_LOGIC_VECTOR (71 DOWNTO 0);
      core_wen1 : IN STD_LOGIC;
      rms_norm_16_div_cmp_z_oreg : OUT STD_LOGIC_VECTOR (39 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL dut_core_wait_dp_inst_rms_norm_16_div_cmp_z : STD_LOGIC_VECTOR (71 DOWNTO
      0);
  SIGNAL dut_core_wait_dp_inst_rms_norm_16_div_cmp_z_oreg : STD_LOGIC_VECTOR (39
      DOWNTO 0);

  COMPONENT dut_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
      for_for_C_2_tr0 : IN STD_LOGIC;
      compute_sqrt_for_C_15_tr0 : IN STD_LOGIC;
      RMS_NORM_LOOP_2_C_4_tr0 : IN STD_LOGIC;
      QUANTIZE_ACTIVATION_LOOP_3_C_2_tr0 : IN STD_LOGIC;
      LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0 : IN STD_LOGIC;
      LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0 : IN STD_LOGIC;
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_63_tr0 : IN STD_LOGIC;
      RESHAPE_2D_TO_3D_LOOP_3_C_0_tr0 : IN STD_LOGIC;
      RESHAPE_2D_TO_3D_LOOP_2_C_0_tr0 : IN STD_LOGIC;
      RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0 : IN STD_LOGIC;
      RESHAPE_2D_TO_3D_LOOP_2_2_C_0_tr0 : IN STD_LOGIC;
      APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0 : IN STD_LOGIC;
      APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0 : IN STD_LOGIC;
      CACHE_UPDATE_LOOP_3_C_1_tr0 : IN STD_LOGIC;
      CACHE_UPDATE_LOOP_2_C_0_tr0 : IN STD_LOGIC;
      CACHE_UPDATE_LOOP_1_C_0_tr0 : IN STD_LOGIC;
      TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0 : IN STD_LOGIC;
      TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0 : IN STD_LOGIC;
      TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0 : IN STD_LOGIC;
      GEMM_3D_FLOAT_LOOP_4_C_3_tr0 : IN STD_LOGIC;
      GEMM_3D_FLOAT_LOOP_3_C_1_tr0 : IN STD_LOGIC;
      GEMM_3D_FLOAT_LOOP_1_C_0_tr0 : IN STD_LOGIC;
      SF_LOOP_3_C_0_tr0 : IN STD_LOGIC;
      SF_LOOP_1_C_0_tr0 : IN STD_LOGIC;
      CM_LOOP_1_C_0_tr0 : IN STD_LOGIC;
      SOFTMAX_LOOP_3_C_0_tr0 : IN STD_LOGIC;
      SOFTMAX_LOOP_4_C_2_tr0 : IN STD_LOGIC;
      SOFTMAX_LOOP_5_C_19_tr0 : IN STD_LOGIC;
      SOFTMAX_LOOP_1_C_1_tr0 : IN STD_LOGIC;
      GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0 : IN STD_LOGIC;
      GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0 : IN STD_LOGIC;
      GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0 : IN STD_LOGIC;
      ATTN_2D_LOOP_3_C_0_tr0 : IN STD_LOGIC;
      ATTN_2D_LOOP_2_C_0_tr0 : IN STD_LOGIC;
      RMS_NORM_LOOP_1_2_C_2_tr0 : IN STD_LOGIC;
      compute_sqrt_1_for_C_15_tr0 : IN STD_LOGIC;
      RMS_NORM_LOOP_2_2_C_4_tr0 : IN STD_LOGIC;
      QUANTIZE_ACTIVATION_LOOP_3_1_C_2_tr0 : IN STD_LOGIC;
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0 : IN STD_LOGIC;
      LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0 : IN STD_LOGIC;
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31_tr0 : IN STD_LOGIC;
      for_1_for_C_1_tr0 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL dut_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL dut_core_core_fsm_inst_compute_sqrt_for_C_15_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_CACHE_UPDATE_LOOP_3_C_1_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_CACHE_UPDATE_LOOP_2_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_3_C_1_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_1_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_SF_LOOP_3_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_SF_LOOP_1_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_CM_LOOP_1_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_SOFTMAX_LOOP_3_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_SOFTMAX_LOOP_4_C_2_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_SOFTMAX_LOOP_5_C_19_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_SOFTMAX_LOOP_1_C_1_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_ATTN_2D_LOOP_3_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_ATTN_2D_LOOP_2_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_compute_sqrt_1_for_C_15_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0 : STD_LOGIC;
  SIGNAL dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_s_1_13_2(input_12 : STD_LOGIC;
  input_11 : STD_LOGIC;
  input_10 : STD_LOGIC;
  input_9 : STD_LOGIC;
  input_8 : STD_LOGIC;
  input_7 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(12 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
      tmp := sel(7);
      result := result or ( input_7 and tmp);
      tmp := sel(8);
      result := result or ( input_8 and tmp);
      tmp := sel(9);
      result := result or ( input_9 and tmp);
      tmp := sel(10);
      result := result or ( input_10 and tmp);
      tmp := sel(11);
      result := result or ( input_11 and tmp);
      tmp := sel(12);
      result := result or ( input_12 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_3_2(input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_4_2(input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_5_2(input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_6_2(input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_7_2(input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_8_2(input_7 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
      tmp := sel(7);
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_9_2(input_8 : STD_LOGIC;
  input_7 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(8 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
      tmp := sel(7);
      result := result or ( input_7 and tmp);
      tmp := sel(8);
      result := result or ( input_8 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_13_3_2(input_2 : STD_LOGIC_VECTOR(12 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(12 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(12 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(12 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(12 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_15_6_2(input_5 : STD_LOGIC_VECTOR(14 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(14 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(14 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(14 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(14 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(14 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(14 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(14 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_16_3_2(input_2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(15 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(15 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_16_4_2(input_3 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(15 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(15 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_16_5_2(input_4 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(15 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(15 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_16_6_2(input_5 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(15 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(15 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_16_7_2(input_6 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(15 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(15 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_16_8_2(input_7 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(15 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(15 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_21_5_2(input_4 : STD_LOGIC_VECTOR(20 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(20 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(20 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(20 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(20 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(20 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(20 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_22_5_2(input_4 : STD_LOGIC_VECTOR(21 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(21 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(21 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(21 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(21 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(21 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(21 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_24_3_2(input_2 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(23 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(23 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_24_4_2(input_3 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(23 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(23 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_24_6_2(input_5 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(23 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(23 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_24_7_2(input_6 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(23 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(23 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_24_8_2(input_7 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(23 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(23 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_24_9_2(input_8 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(8 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(23 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(23 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_2_6_2(input_5 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_2_7_2(input_6 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_34_7_2(input_6 : STD_LOGIC_VECTOR(33 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(33 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(33 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(33 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(33 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(33 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(33 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(33 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(33 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_38_5_2(input_4 : STD_LOGIC_VECTOR(37 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(37 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(37 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(37 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(37 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(37 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(37 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_39_10_2(input_9 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(9 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(38 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(38 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_39_13_2(input_12 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(12 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(38 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(38 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_39_3_2(input_2 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(38 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(38 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_39_5_2(input_4 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(38 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(38 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_39_8_2(input_7 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(38 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(38 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_3_2(input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_4_2(input_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_5_2(input_4 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_6_2(input_5 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_40_10_2(input_9 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(9 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(39 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(39 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_40_11_2(input_10 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(10 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(39 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(39 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_40_3_2(input_2 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(39 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(39 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_40_6_2(input_5 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(39 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(39 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_40_7_2(input_6 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(39 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(39 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_40_8_2(input_7 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(39 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(39 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_40_9_2(input_8 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(8 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(39 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(39 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_5_2(input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_6_2(input_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_5_6_2(input_5 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_5_7_2(input_6 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_6_2(input_5 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_7_7_2(input_6 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_8_3_2(input_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_8_4_2(input_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_8_6_2(input_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_8_7_2(input_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_8_8_2(input_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_8_9_2(input_8 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(8 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_16_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_7 : STD_LOGIC;
  input_8 : STD_LOGIC;
  input_9 : STD_LOGIC;
  input_10 : STD_LOGIC;
  input_11 : STD_LOGIC;
  input_12 : STD_LOGIC;
  input_13 : STD_LOGIC;
  input_14 : STD_LOGIC;
  input_15 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN "1001" =>
          result := input_9;
        WHEN "1010" =>
          result := input_10;
        WHEN "1011" =>
          result := input_11;
        WHEN "1100" =>
          result := input_12;
        WHEN "1101" =>
          result := input_13;
        WHEN "1110" =>
          result := input_14;
        WHEN others =>
          result := input_15;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_s_1_4_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_3 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(1 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN "00" =>
          result := input_0;
        WHEN "01" =>
          result := input_1;
        WHEN "10" =>
          result := input_2;
        WHEN others =>
          result := input_3;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_s_1_8_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_7 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN "000" =>
          result := input_0;
        WHEN "001" =>
          result := input_1;
        WHEN "010" =>
          result := input_2;
        WHEN "011" =>
          result := input_3;
        WHEN "100" =>
          result := input_4;
        WHEN "101" =>
          result := input_5;
        WHEN "110" =>
          result := input_6;
        WHEN others =>
          result := input_7;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_12_16_2(input_0 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(11 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN "1001" =>
          result := input_9;
        WHEN "1010" =>
          result := input_10;
        WHEN "1011" =>
          result := input_11;
        WHEN "1100" =>
          result := input_12;
        WHEN "1101" =>
          result := input_13;
        WHEN "1110" =>
          result := input_14;
        WHEN others =>
          result := input_15;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_13_2_2(input_0 : STD_LOGIC_VECTOR(12 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(12 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(12 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_14_16_2(input_0 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(13 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN "1001" =>
          result := input_9;
        WHEN "1010" =>
          result := input_10;
        WHEN "1011" =>
          result := input_11;
        WHEN "1100" =>
          result := input_12;
        WHEN "1101" =>
          result := input_13;
        WHEN "1110" =>
          result := input_14;
        WHEN others =>
          result := input_15;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_14_2_2(input_0 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(13 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_16_16_2(input_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(15 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN "1001" =>
          result := input_9;
        WHEN "1010" =>
          result := input_10;
        WHEN "1011" =>
          result := input_11;
        WHEN "1100" =>
          result := input_12;
        WHEN "1101" =>
          result := input_13;
        WHEN "1110" =>
          result := input_14;
        WHEN others =>
          result := input_15;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_16_2_2(input_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(15 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_23_16_2(input_0 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(22 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(22 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN "1001" =>
          result := input_9;
        WHEN "1010" =>
          result := input_10;
        WHEN "1011" =>
          result := input_11;
        WHEN "1100" =>
          result := input_12;
        WHEN "1101" =>
          result := input_13;
        WHEN "1110" =>
          result := input_14;
        WHEN others =>
          result := input_15;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_24_16_2(input_0 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(23 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN "1001" =>
          result := input_9;
        WHEN "1010" =>
          result := input_10;
        WHEN "1011" =>
          result := input_11;
        WHEN "1100" =>
          result := input_12;
        WHEN "1101" =>
          result := input_13;
        WHEN "1110" =>
          result := input_14;
        WHEN others =>
          result := input_15;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_24_2_2(input_0 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(23 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_24_8_2(input_0 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(23 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(23 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "000" =>
          result := input_0;
        WHEN "001" =>
          result := input_1;
        WHEN "010" =>
          result := input_2;
        WHEN "011" =>
          result := input_3;
        WHEN "100" =>
          result := input_4;
        WHEN "101" =>
          result := input_5;
        WHEN "110" =>
          result := input_6;
        WHEN others =>
          result := input_7;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_2_2_2(input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_2_4_2(input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(1 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "00" =>
          result := input_0;
        WHEN "01" =>
          result := input_1;
        WHEN "10" =>
          result := input_2;
        WHEN others =>
          result := input_3;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_34_2_2(input_0 : STD_LOGIC_VECTOR(33 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(33 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(33 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_35_2_2(input_0 : STD_LOGIC_VECTOR(34 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(34 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(34 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_39_16_2(input_0 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(38 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN "1001" =>
          result := input_9;
        WHEN "1010" =>
          result := input_10;
        WHEN "1011" =>
          result := input_11;
        WHEN "1100" =>
          result := input_12;
        WHEN "1101" =>
          result := input_13;
        WHEN "1110" =>
          result := input_14;
        WHEN others =>
          result := input_15;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_39_2_2(input_0 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(38 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(38 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_3_16_2(input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN "1001" =>
          result := input_9;
        WHEN "1010" =>
          result := input_10;
        WHEN "1011" =>
          result := input_11;
        WHEN "1100" =>
          result := input_12;
        WHEN "1101" =>
          result := input_13;
        WHEN "1110" =>
          result := input_14;
        WHEN others =>
          result := input_15;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_3_2_2(input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_3_8_2(input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "000" =>
          result := input_0;
        WHEN "001" =>
          result := input_1;
        WHEN "010" =>
          result := input_2;
        WHEN "011" =>
          result := input_3;
        WHEN "100" =>
          result := input_4;
        WHEN "101" =>
          result := input_5;
        WHEN "110" =>
          result := input_6;
        WHEN others =>
          result := input_7;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_40_12_2(input_0 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(39 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN "1001" =>
          result := input_9;
        WHEN "1010" =>
          result := input_10;
        WHEN others =>
          result := input_11;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_40_15_2(input_0 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(39 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN "1001" =>
          result := input_9;
        WHEN "1010" =>
          result := input_10;
        WHEN "1011" =>
          result := input_11;
        WHEN "1100" =>
          result := input_12;
        WHEN "1101" =>
          result := input_13;
        WHEN others =>
          result := input_14;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_40_16_2(input_0 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(39 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN "1001" =>
          result := input_9;
        WHEN "1010" =>
          result := input_10;
        WHEN "1011" =>
          result := input_11;
        WHEN "1100" =>
          result := input_12;
        WHEN "1101" =>
          result := input_13;
        WHEN "1110" =>
          result := input_14;
        WHEN others =>
          result := input_15;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_40_2_2(input_0 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(39 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_40_4_2(input_0 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(39 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(1 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(39 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "00" =>
          result := input_0;
        WHEN "01" =>
          result := input_1;
        WHEN "10" =>
          result := input_2;
        WHEN others =>
          result := input_3;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_4_2_2(input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_53_2_2(input_0 : STD_LOGIC_VECTOR(52 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(52 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(52 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_7_2_2(input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_8_16_2(input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN "1001" =>
          result := input_9;
        WHEN "1010" =>
          result := input_10;
        WHEN "1011" =>
          result := input_11;
        WHEN "1100" =>
          result := input_12;
        WHEN "1101" =>
          result := input_13;
        WHEN "1110" =>
          result := input_14;
        WHEN others =>
          result := input_15;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_8_2_2(input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_8_8_2(input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "000" =>
          result := input_0;
        WHEN "001" =>
          result := input_1;
        WHEN "010" =>
          result := input_2;
        WHEN "011" =>
          result := input_3;
        WHEN "100" =>
          result := input_4;
        WHEN "101" =>
          result := input_5;
        WHEN "110" =>
          result := input_6;
        WHEN others =>
          result := input_7;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_9_16_2(input_0 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(8 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN "1001" =>
          result := input_9;
        WHEN "1010" =>
          result := input_10;
        WHEN "1011" =>
          result := input_11;
        WHEN "1100" =>
          result := input_12;
        WHEN "1101" =>
          result := input_13;
        WHEN "1110" =>
          result := input_14;
        WHEN others =>
          result := input_15;
      END CASE;
    RETURN result;
  END;

BEGIN
  SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp : work.mgc_comps.mgc_div
    GENERIC MAP(
      width_a => 56,
      width_b => 40,
      signd => 1
      )
    PORT MAP(
      a => SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a,
      b => SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b,
      z => SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z_1
    );
  SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a <= SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_55
      & SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_54_16 & STD_LOGIC_VECTOR'( "0000000000000000");
  SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b <= SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_39
      & SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_38_0;
  SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z <= SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z_1;

  LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp : work.mgc_comps.mgc_div
    GENERIC MAP(
      width_a => 72,
      width_b => 60,
      signd => 1
      )
    PORT MAP(
      a => LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a,
      b => LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b,
      z => LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z_1
    );
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a <= LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_71_48
      & LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_47_40
      & LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_39
      & LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_38
      & LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_37
      & LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_36
      & LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_35
      & LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_34
      & LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_33
      & LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_32
      & STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b <= LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_59_39
      & LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_38_0;
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z <= LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z_1;

  operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp : work.mgc_comps.mgc_div
    GENERIC MAP(
      width_a => 40,
      width_b => 40,
      signd => 1
      )
    PORT MAP(
      a => operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a,
      b => operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b,
      z => operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_1
    );
  operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a <= STD_LOGIC_VECTOR(UNSIGNED'( "0")
      & UNSIGNED(CONV_SIGNED(SIGNED(reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd
      & STD_LOGIC_VECTOR'( "000000000000000") & reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd_1
      & STD_LOGIC_VECTOR'( "0000000000000000")),39)));
  operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b <= operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_39
      & operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_38_35 & operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_34
      & operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_33_0;
  operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z <= operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_1;

  CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_rg : work.dutmgc_rom_33_32_20_1_pkg.dutmgc_rom_33_32_20_1
    PORT MAP(
      addr => CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_rg_addr,
      data_out => CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_rg_data_out
    );
  CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_rg_addr <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd,
      1), 1), 2) + UNSIGNED'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1),
      2)) & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1;
  CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_sdt <= CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_rg_data_out;

  LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_rg : work.dutmgc_rom_34_64_8_1_pkg.dutmgc_rom_34_64_8_1
    PORT MAP(
      addr => LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_rg_addr,
      data_out => LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_rg_data_out
    );
  LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_rg_addr
      <= reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2;
  LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_itm <= LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_rg_data_out;

  LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_rg : work.dutmgc_rom_35_64_8_1_pkg.dutmgc_rom_35_64_8_1
    PORT MAP(
      addr => LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_rg_addr,
      data_out => LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_rg_data_out
    );
  LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_rg_addr
      <= reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2;
  LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_itm <= LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_rg_data_out;

  APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_rg : work.dutmgc_rom_36_960_15_1_pkg.dutmgc_rom_36_960_15_1
    PORT MAP(
      addr => APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_rg_addr,
      data_out => APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_rg_data_out
    );
  APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_rg_addr <= STD_LOGIC_VECTOR'(
      "00110000") & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1;
  APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_itm <= APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_rg_data_out;

  APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_rg : work.dutmgc_rom_37_960_13_1_pkg.dutmgc_rom_37_960_13_1
    PORT MAP(
      addr => APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_rg_addr,
      data_out => APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_rg_data_out
    );
  APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_rg_addr <= STD_LOGIC_VECTOR'(
      "00110000") & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1;
  APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm <= APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_rg_data_out;

  LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_rg : work.dutmgc_rom_38_64_8_1_pkg.dutmgc_rom_38_64_8_1
    PORT MAP(
      addr => LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_rg_addr,
      data_out => LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_rg_data_out
    );
  LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_rg_addr
      <= reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm <= LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_rg_data_out;

  LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_rg : work.dutmgc_rom_39_64_8_1_pkg.dutmgc_rom_39_64_8_1
    PORT MAP(
      addr => LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_rg_addr,
      data_out => LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_rg_data_out
    );
  LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_rg_addr <=
      reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 &
      reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1;
  LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm <= LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_rg_data_out;

  CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_rg : work.dutmgc_rom_40_32_19_1_pkg.dutmgc_rom_40_32_19_1
    PORT MAP(
      addr => CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_rg_addr,
      data_out => CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_rg_data_out
    );
  CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_rg_addr <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(1),
      1), 1), 2) + UNSIGNED'( reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1),
      2)) & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0)) & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_itm <= CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_rg_data_out;

  dut_core_strm_in_rsci_inst : dut_core_strm_in_rsci
    PORT MAP(
      strm_in_rsc_dat => dut_core_strm_in_rsci_inst_strm_in_rsc_dat,
      strm_in_rsc_vld => strm_in_rsc_vld,
      strm_in_rsc_rdy => strm_in_rsc_rdy,
      strm_in_rsci_oswt => reg_strm_in_rsci_iswt0_cse,
      strm_in_rsci_wen_comp => strm_in_rsci_wen_comp,
      strm_in_rsci_idat_mxwt => dut_core_strm_in_rsci_inst_strm_in_rsci_idat_mxwt
    );
  dut_core_strm_in_rsci_inst_strm_in_rsc_dat <= strm_in_rsc_dat;
  strm_in_rsci_idat_mxwt <= dut_core_strm_in_rsci_inst_strm_in_rsci_idat_mxwt;

  dut_core_strm_out_rsci_inst : dut_core_strm_out_rsci
    PORT MAP(
      strm_out_rsc_dat => dut_core_strm_out_rsci_inst_strm_out_rsc_dat,
      strm_out_rsc_vld => strm_out_rsc_vld,
      strm_out_rsc_rdy => strm_out_rsc_rdy,
      strm_out_rsci_oswt => reg_strm_out_rsci_iswt0_cse,
      strm_out_rsci_wen_comp => strm_out_rsci_wen_comp,
      strm_out_rsci_idat => dut_core_strm_out_rsci_inst_strm_out_rsci_idat
    );
  strm_out_rsc_dat <= dut_core_strm_out_rsci_inst_strm_out_rsc_dat;
  dut_core_strm_out_rsci_inst_strm_out_rsci_idat <= strm_out_rsci_idat_31_18 & strm_out_rsci_idat_17_10
      & strm_out_rsci_idat_9 & strm_out_rsci_idat_8 & strm_out_rsci_idat_7 & strm_out_rsci_idat_6
      & strm_out_rsci_idat_5 & strm_out_rsci_idat_4 & strm_out_rsci_idat_3 & strm_out_rsci_idat_2
      & STD_LOGIC_VECTOR'( "00");

  dut_core_staller_inst : dut_core_staller
    PORT MAP(
      en => en,
      core_wen1 => core_wen1,
      strm_in_rsci_wen_comp => strm_in_rsci_wen_comp,
      strm_out_rsci_wen_comp => strm_out_rsci_wen_comp,
      attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 => attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
    );
  dut_core_wait_dp_inst : dut_core_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      rms_norm_16_div_cmp_z => dut_core_wait_dp_inst_rms_norm_16_div_cmp_z,
      core_wen1 => core_wen1,
      rms_norm_16_div_cmp_z_oreg => dut_core_wait_dp_inst_rms_norm_16_div_cmp_z_oreg
    );
  dut_core_wait_dp_inst_rms_norm_16_div_cmp_z <= rms_norm_16_div_cmp_z;
  rms_norm_16_div_cmp_z_oreg <= dut_core_wait_dp_inst_rms_norm_16_div_cmp_z_oreg;

  dut_core_core_fsm_inst : dut_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 => attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1,
      fsm_output => dut_core_core_fsm_inst_fsm_output,
      for_for_C_2_tr0 => for_for_and_tmp,
      compute_sqrt_for_C_15_tr0 => dut_core_core_fsm_inst_compute_sqrt_for_C_15_tr0,
      RMS_NORM_LOOP_2_C_4_tr0 => and_37_cse,
      QUANTIZE_ACTIVATION_LOOP_3_C_2_tr0 => LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4,
      LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0 => dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0,
      LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0 => dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_63_tr0 => reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1,
      RESHAPE_2D_TO_3D_LOOP_3_C_0_tr0 => CACHE_UPDATE_LOOP_1_and_tmp,
      RESHAPE_2D_TO_3D_LOOP_2_C_0_tr0 => RESHAPE_2D_TO_3D_LOOP_2_2_and_cse,
      RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0 => dut_core_core_fsm_inst_RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0,
      RESHAPE_2D_TO_3D_LOOP_2_2_C_0_tr0 => RESHAPE_2D_TO_3D_LOOP_2_2_and_cse,
      APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0 => dut_core_core_fsm_inst_APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0,
      APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0 => dut_core_core_fsm_inst_APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0,
      CACHE_UPDATE_LOOP_3_C_1_tr0 => dut_core_core_fsm_inst_CACHE_UPDATE_LOOP_3_C_1_tr0,
      CACHE_UPDATE_LOOP_2_C_0_tr0 => dut_core_core_fsm_inst_CACHE_UPDATE_LOOP_2_C_0_tr0,
      CACHE_UPDATE_LOOP_1_C_0_tr0 => CACHE_UPDATE_LOOP_1_and_tmp,
      TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0 => dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0,
      TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0 => dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0,
      TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0 => dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0,
      GEMM_3D_FLOAT_LOOP_4_C_3_tr0 => reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1,
      GEMM_3D_FLOAT_LOOP_3_C_1_tr0 => dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_3_C_1_tr0,
      GEMM_3D_FLOAT_LOOP_1_C_0_tr0 => dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_1_C_0_tr0,
      SF_LOOP_3_C_0_tr0 => dut_core_core_fsm_inst_SF_LOOP_3_C_0_tr0,
      SF_LOOP_1_C_0_tr0 => dut_core_core_fsm_inst_SF_LOOP_1_C_0_tr0,
      CM_LOOP_1_C_0_tr0 => dut_core_core_fsm_inst_CM_LOOP_1_C_0_tr0,
      SOFTMAX_LOOP_3_C_0_tr0 => dut_core_core_fsm_inst_SOFTMAX_LOOP_3_C_0_tr0,
      SOFTMAX_LOOP_4_C_2_tr0 => dut_core_core_fsm_inst_SOFTMAX_LOOP_4_C_2_tr0,
      SOFTMAX_LOOP_5_C_19_tr0 => dut_core_core_fsm_inst_SOFTMAX_LOOP_5_C_19_tr0,
      SOFTMAX_LOOP_1_C_1_tr0 => dut_core_core_fsm_inst_SOFTMAX_LOOP_1_C_1_tr0,
      GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0 => dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0,
      GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0 => dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0,
      GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0 => dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0,
      ATTN_2D_LOOP_3_C_0_tr0 => dut_core_core_fsm_inst_ATTN_2D_LOOP_3_C_0_tr0,
      ATTN_2D_LOOP_2_C_0_tr0 => dut_core_core_fsm_inst_ATTN_2D_LOOP_2_C_0_tr0,
      RMS_NORM_LOOP_1_2_C_2_tr0 => LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4,
      compute_sqrt_1_for_C_15_tr0 => dut_core_core_fsm_inst_compute_sqrt_1_for_C_15_tr0,
      RMS_NORM_LOOP_2_2_C_4_tr0 => and_37_cse,
      QUANTIZE_ACTIVATION_LOOP_3_1_C_2_tr0 => LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4,
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0 => dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0,
      LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0 => dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0,
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31_tr0 => LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4,
      for_1_for_C_1_tr0 => LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4
    );
  fsm_output <= dut_core_core_fsm_inst_fsm_output;
  dut_core_core_fsm_inst_compute_sqrt_for_C_15_tr0 <= NOT reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0 <= (LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_2(2))
      AND (z_out_5(2)) AND (z_out_3(2));
  dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0 <= (z_out_3(2)) AND
      (z_out_4(2)) AND (z_out_5(2));
  dut_core_core_fsm_inst_RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0 <= (reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      OR reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1) AND (z_out_3(2));
  dut_core_core_fsm_inst_APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0 <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1);
  dut_core_core_fsm_inst_APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0 <= z_out_4(2);
  dut_core_core_fsm_inst_CACHE_UPDATE_LOOP_3_C_1_tr0 <= reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1
      AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1));
  dut_core_core_fsm_inst_CACHE_UPDATE_LOOP_2_C_0_tr0 <= NOT(CACHE_UPDATE_LOOP_2_acc_2_itm_2_1
      OR CACHE_UPDATE_LOOP_2_1_acc_2_itm_2_1);
  dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0 <= TRANSPOSE_LAST_TWO_DIMS_LOOP_3_k_2_0_sva_1(2);
  dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0 <= NOT CACHE_UPDATE_LOOP_2_1_acc_2_itm_2_1;
  dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0 <= z_out_5(2);
  dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_3_C_1_tr0 <= NOT CACHE_UPDATE_LOOP_2_1_acc_2_itm_2_1;
  dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_1_C_0_tr0 <= z_out_5(2);
  dut_core_core_fsm_inst_SF_LOOP_3_C_0_tr0 <= NOT CACHE_UPDATE_LOOP_2_1_acc_2_itm_2_1;
  dut_core_core_fsm_inst_SF_LOOP_1_C_0_tr0 <= z_out_5(2);
  dut_core_core_fsm_inst_CM_LOOP_1_C_0_tr0 <= z_out_3(2);
  dut_core_core_fsm_inst_SOFTMAX_LOOP_3_C_0_tr0 <= NOT reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  dut_core_core_fsm_inst_SOFTMAX_LOOP_4_C_2_tr0 <= NOT reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  dut_core_core_fsm_inst_SOFTMAX_LOOP_5_C_19_tr0 <= NOT reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  dut_core_core_fsm_inst_SOFTMAX_LOOP_1_C_1_tr0 <= z_out_5(2);
  dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0 <= NOT reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0 <= z_out_4(2);
  dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0 <= z_out_5(2);
  dut_core_core_fsm_inst_ATTN_2D_LOOP_3_C_0_tr0 <= z_out_5(2);
  dut_core_core_fsm_inst_ATTN_2D_LOOP_2_C_0_tr0 <= z_out_4(2);
  dut_core_core_fsm_inst_compute_sqrt_1_for_C_15_tr0 <= NOT reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0 <= z_out_5(2);
  dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0 <= z_out_4(2);

  attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1;
  for_1_for_and_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT(or_dcpl_961
      OR (NOT((fsm_output(5)) AND (fsm_output(3)))) OR or_1984_cse));
  attention_2_1_16_16_4_4_attn_output_and_4_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND and_dcpl_187;
  nand_302_cse <= NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd AND GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva);
  nand_303_tmp <= NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd AND GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva);
  attention_2_1_16_16_4_4_attn_output_and_14_cse <= nand_303_tmp AND and_dcpl_187;
  attention_2_1_16_16_4_4_attn_output_and_13_cse <= (NOT nand_303_tmp) AND and_dcpl_187;
  nand_304_tmp <= NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd AND GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva);
  attention_2_1_16_16_4_4_attn_output_and_16_cse <= nand_304_tmp AND and_dcpl_187;
  attention_2_1_16_16_4_4_attn_output_and_15_cse <= (NOT nand_304_tmp) AND and_dcpl_187;
  nand_305_tmp <= NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd AND GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva);
  attention_2_1_16_16_4_4_attn_output_and_18_cse <= nand_305_tmp AND and_dcpl_187;
  attention_2_1_16_16_4_4_attn_output_and_17_cse <= (NOT nand_305_tmp) AND and_dcpl_187;
  and_1481_nl <= (((fsm_output(2)) AND (fsm_output(6))) OR (fsm_output(7))) AND (fsm_output(8));
  mux_775_nl <= MUX_s_1_2_2(and_1481_nl, mux_tmp_363, fsm_output(5));
  or_1677_nl <= (z_out_5(2)) OR (NOT (fsm_output(5))) OR (fsm_output(2));
  mux_774_nl <= MUX_s_1_2_2(mux_tmp_363, nor_tmp_117, or_1677_nl);
  mux_776_nl <= MUX_s_1_2_2(mux_775_nl, mux_774_nl, fsm_output(3));
  or_1676_nl <= (fsm_output(3)) OR (NOT (fsm_output(5))) OR (fsm_output(2));
  mux_773_nl <= MUX_s_1_2_2(mux_tmp_363, nor_tmp_117, or_1676_nl);
  mux_777_nl <= MUX_s_1_2_2(mux_776_nl, mux_773_nl, or_1732_cse);
  mux_778_nl <= MUX_s_1_2_2(mux_777_nl, nor_tmp_117, fsm_output(4));
  attention_2_1_16_16_4_4_attn_weights_and_36_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND mux_778_nl;
  attention_2_1_16_16_4_4_q_embed_and_5_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND and_dcpl_204;
  attention_2_1_16_16_4_4_q_embed_and_23_cse <= (NOT or_dcpl_991) AND and_dcpl_204;
  attention_2_1_16_16_4_4_q_embed_and_24_cse <= or_dcpl_991 AND and_dcpl_204;
  attention_2_1_16_16_4_4_q_embed_mux_7_cse <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_q_embed_2_0_3_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1, attention_2_1_16_16_4_4_q_embed_2_0_3_lpi_3,
      STD_LOGIC_VECTOR'( (NOT and_dcpl_204) & attention_2_1_16_16_4_4_q_embed_and_23_cse
      & attention_2_1_16_16_4_4_q_embed_and_24_cse));
  attention_2_1_16_16_4_4_q_embed_and_25_cse <= (NOT or_dcpl_995) AND and_dcpl_204;
  attention_2_1_16_16_4_4_q_embed_and_26_cse <= or_dcpl_995 AND and_dcpl_204;
  attention_2_1_16_16_4_4_q_embed_mux_9_cse <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_q_embed_3_0_0_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1, attention_2_1_16_16_4_4_q_embed_3_0_0_lpi_3,
      STD_LOGIC_VECTOR'( (NOT and_dcpl_204) & attention_2_1_16_16_4_4_q_embed_and_25_cse
      & attention_2_1_16_16_4_4_q_embed_and_26_cse));
  attention_2_1_16_16_4_4_q_embed_and_27_cse <= (NOT or_dcpl_997) AND and_dcpl_204;
  attention_2_1_16_16_4_4_q_embed_and_28_cse <= or_dcpl_997 AND and_dcpl_204;
  attention_2_1_16_16_4_4_q_embed_mux_11_cse <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_q_embed_3_0_1_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1, attention_2_1_16_16_4_4_q_embed_3_0_1_lpi_3,
      STD_LOGIC_VECTOR'( (NOT and_dcpl_204) & attention_2_1_16_16_4_4_q_embed_and_27_cse
      & attention_2_1_16_16_4_4_q_embed_and_28_cse));
  attention_2_1_16_16_4_4_q_embed_and_29_cse <= (NOT or_dcpl_999) AND and_dcpl_204;
  attention_2_1_16_16_4_4_q_embed_and_30_cse <= or_dcpl_999 AND and_dcpl_204;
  attention_2_1_16_16_4_4_q_embed_mux_13_cse <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_q_embed_3_0_2_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1, attention_2_1_16_16_4_4_q_embed_3_0_2_lpi_3,
      STD_LOGIC_VECTOR'( (NOT and_dcpl_204) & attention_2_1_16_16_4_4_q_embed_and_29_cse
      & attention_2_1_16_16_4_4_q_embed_and_30_cse));
  attention_2_1_16_16_4_4_q_embed_and_31_nl <= (NOT or_dcpl_1000) AND and_dcpl_204;
  attention_2_1_16_16_4_4_q_embed_and_32_nl <= or_dcpl_1000 AND and_dcpl_204;
  attention_2_1_16_16_4_4_q_embed_mux_14_cse <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_q_embed_3_0_3_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1, attention_2_1_16_16_4_4_q_embed_3_0_3_lpi_3,
      STD_LOGIC_VECTOR'( (NOT and_dcpl_204) & attention_2_1_16_16_4_4_q_embed_and_31_nl
      & attention_2_1_16_16_4_4_q_embed_and_32_nl));
  attention_2_1_16_16_4_4_v_proj_and_2_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND and_dcpl_207;
  nor_728_nl <= NOT((fsm_output(4)) OR (fsm_output(7)));
  mux_781_nl <= MUX_s_1_2_2(nor_728_nl, (fsm_output(7)), fsm_output(6));
  mux_782_nl <= MUX_s_1_2_2(mux_781_nl, and_dcpl_148, fsm_output(2));
  mux_783_nl <= MUX_s_1_2_2(mux_782_nl, nor_tmp_261, fsm_output(1));
  and_1383_nl <= (fsm_output(4)) AND (fsm_output(7));
  mux_779_nl <= MUX_s_1_2_2(and_dcpl_148, and_1383_nl, fsm_output(2));
  mux_780_nl <= MUX_s_1_2_2(nor_tmp_261, mux_779_nl, fsm_output(1));
  mux_784_nl <= MUX_s_1_2_2(mux_783_nl, mux_780_nl, fsm_output(0));
  and_1485_nl <= or_1879_cse AND (fsm_output(7));
  mux_785_nl <= MUX_s_1_2_2(mux_784_nl, and_1485_nl, fsm_output(3));
  mux_786_nl <= MUX_s_1_2_2(mux_785_nl, (fsm_output(7)), fsm_output(5));
  apply_rotary_pos_emb_1_4_4_rotated_q_and_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (mux_786_nl OR (fsm_output(8)));
  apply_rotary_pos_emb_1_4_4_rotated_q_or_11_cse <= (and_dcpl_186 AND and_dcpl_209)
      OR ((NOT RESHAPE_2D_TO_3D_LOOP_2_2_and_cse) AND and_dcpl_213);
  apply_rotary_pos_emb_1_4_4_rotated_q_or_12_cse <= (RESHAPE_2D_TO_3D_LOOP_2_2_and_cse
      AND and_dcpl_213) OR and_dcpl_216;
  or_1732_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"));
  mux_792_cse <= MUX_s_1_2_2((fsm_output(7)), (NOT (fsm_output(7))), fsm_output(6));
  attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1 <= MUX_v_24_16_2(attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_3_39_16, apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_39_16,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16, attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_3_39_16, attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_3_39_16, attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_3_39_16, attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_3_39_16, attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_3_39_16, attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_3_39_16, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  attention_2_1_16_16_4_4_q_proj_and_23_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND and_dcpl_240;
  RESHAPE_2D_TO_3D_LOOP_3_1_mux_13_cse <= MUX_v_8_2_2((z_out_1(15 DOWNTO 8)), LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8,
      or_dcpl_1011);
  RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_7 <= MUX_s_1_2_2((z_out_1(7)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd,
      or_dcpl_1011);
  RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_6 <= MUX_s_1_2_2((z_out_1(6)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1,
      or_dcpl_1011);
  RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_5 <= MUX_s_1_2_2((z_out_1(5)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2,
      or_dcpl_1011);
  RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_4 <= MUX_s_1_2_2((z_out_1(4)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3,
      or_dcpl_1011);
  RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_3 <= MUX_s_1_2_2((z_out_1(3)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4,
      or_dcpl_1011);
  RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_2 <= MUX_s_1_2_2((z_out_1(2)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5,
      or_dcpl_1011);
  RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_1 <= MUX_s_1_2_2((z_out_1(1)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6,
      or_dcpl_1011);
  RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_0 <= MUX_s_1_2_2((z_out_1(0)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7,
      or_dcpl_1011);
  and_274_nl <= or_1732_cse AND mux_tmp_121;
  mux_801_nl <= MUX_s_1_2_2(and_274_nl, nor_tmp_28, or_2699_cse);
  nor_271_nl <= NOT(and_37_cse OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")));
  mux_799_nl <= MUX_s_1_2_2(nor_tmp_28, mux_tmp_121, nor_271_nl);
  mux_800_nl <= MUX_s_1_2_2(nor_tmp_28, mux_799_nl, and_1762_cse);
  mux_802_nl <= MUX_s_1_2_2(mux_801_nl, mux_800_nl, fsm_output(3));
  mux_803_nl <= MUX_s_1_2_2(mux_802_nl, nor_tmp_28, fsm_output(2));
  mux_804_nl <= MUX_s_1_2_2(mux_803_nl, (fsm_output(8)), fsm_output(7));
  input_and_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND mux_804_nl;
  and_1555_cse <= (fsm_output(0)) AND (fsm_output(2));
  or_1769_cse <= (NOT (fsm_output(5))) OR (fsm_output(8));
  or_1770_cse <= (fsm_output(5)) OR (NOT (fsm_output(8)));
  and_1559_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  mux_806_cse <= MUX_s_1_2_2((NOT (fsm_output(7))), (fsm_output(7)), fsm_output(6));
  nor_973_cse <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  or_270_cse <= (NOT (fsm_output(2))) OR (fsm_output(4));
  or_1767_cse <= (NOT (fsm_output(7))) OR (fsm_output(5)) OR (fsm_output(8));
  or_1772_cse <= (fsm_output(4)) OR (fsm_output(7)) OR (fsm_output(5)) OR (fsm_output(8));
  or_1775_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(5)) OR (fsm_output(8));
  or_1774_nl <= (fsm_output(1)) OR and_1555_cse OR (fsm_output(7)) OR (fsm_output(5))
      OR (fsm_output(8));
  mux_814_nl <= MUX_s_1_2_2(or_1775_nl, or_1774_nl, fsm_output(4));
  mux_815_nl <= MUX_s_1_2_2(mux_814_nl, or_1772_cse, fsm_output(3));
  mux_811_nl <= MUX_s_1_2_2(or_1770_cse, or_1769_cse, fsm_output(7));
  or_1771_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR
      mux_811_nl;
  mux_812_nl <= MUX_s_1_2_2(or_1771_nl, or_1767_cse, fsm_output(4));
  nand_41_nl <= NOT((fsm_output(4)) AND (NOT(and_1559_cse OR (NOT (fsm_output(7)))
      OR (fsm_output(5)) OR (fsm_output(8)))));
  mux_813_nl <= MUX_s_1_2_2(mux_812_nl, nand_41_nl, fsm_output(3));
  mux_816_ssc <= MUX_s_1_2_2(mux_815_nl, mux_813_nl, fsm_output(6));
  and_303_ssc <= (NOT mux_tmp_836) AND and_dcpl_270;
  compute_sqrt_guess_or_1_ssc <= ((NOT and_dcpl_290) AND and_dcpl_272 AND nor_777_cse
      AND and_dcpl_209) OR ((NOT and_dcpl_292) AND and_dcpl_226 AND (NOT (fsm_output(1)))
      AND ((fsm_output(4)) XOR (fsm_output(5))) AND (NOT((fsm_output(0)) OR (fsm_output(3))))
      AND and_dcpl_148);
  mux_838_nl <= MUX_s_1_2_2(or_3185_cse, (NOT and_1559_cse), fsm_output(3));
  and_315_ssc <= mux_838_nl AND (NOT (fsm_output(8))) AND and_dcpl_279 AND and_dcpl_148;
  or_1803_nl <= (fsm_output(1)) OR (NOT (fsm_output(4))) OR (fsm_output(7)) OR (fsm_output(5))
      OR (fsm_output(8));
  mux_848_nl <= MUX_s_1_2_2(or_1772_cse, mux_tmp_841, fsm_output(1));
  mux_849_nl <= MUX_s_1_2_2(or_1803_nl, mux_848_nl, fsm_output(3));
  mux_845_nl <= MUX_s_1_2_2((fsm_output(5)), or_1769_cse, fsm_output(7));
  or_1802_nl <= (fsm_output(4)) OR mux_845_nl;
  mux_846_nl <= MUX_s_1_2_2(or_1802_nl, mux_tmp_839, or_1732_cse);
  or_1799_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(7))) OR (fsm_output(5))
      OR (fsm_output(8));
  mux_847_nl <= MUX_s_1_2_2(mux_846_nl, or_1799_nl, fsm_output(3));
  mux_850_nl <= MUX_s_1_2_2(mux_849_nl, mux_847_nl, fsm_output(6));
  or_1798_nl <= (NOT (fsm_output(4))) OR (fsm_output(7)) OR (fsm_output(5)) OR (fsm_output(8));
  mux_842_nl <= MUX_s_1_2_2(or_1798_nl, or_1772_cse, or_1732_cse);
  mux_843_nl <= MUX_s_1_2_2(mux_842_nl, mux_tmp_841, fsm_output(3));
  or_1792_nl <= (fsm_output(1)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(7)))
      OR (fsm_output(5)) OR (fsm_output(8));
  mux_840_nl <= MUX_s_1_2_2(mux_tmp_839, or_1792_nl, fsm_output(3));
  mux_844_nl <= MUX_s_1_2_2(mux_843_nl, mux_840_nl, fsm_output(6));
  mux_851_ssc <= MUX_s_1_2_2(mux_850_nl, mux_844_nl, fsm_output(2));
  nor_977_nl <= NOT((fsm_output(6)) OR mux_tmp_836);
  and_1561_nl <= (NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))))
      AND (fsm_output(4));
  mux_852_nl <= MUX_s_1_2_2(nor_tmp_285, and_1561_nl, fsm_output(3));
  and_1562_nl <= (fsm_output(6)) AND mux_852_nl;
  mux_853_nl <= MUX_s_1_2_2(nor_977_nl, and_1562_nl, fsm_output(7));
  and_321_ssc <= mux_853_nl AND and_dcpl_1;
  and_1474_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  mux_854_nl <= MUX_s_1_2_2(and_1762_cse, (NOT or_tmp_755), fsm_output(6));
  and_329_ssc <= mux_854_nl AND and_dcpl_295;
  and_334_ssc <= (NOT((NOT(nand_197_cse AND CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("00"))))
      AND (fsm_output(4)))) AND and_dcpl_298;
  and_336_ssc <= and_dcpl_206 AND and_dcpl_302;
  or_1812_nl <= (fsm_output(5)) OR (fsm_output(4)) OR (NOT (fsm_output(8)));
  mux_855_nl <= MUX_s_1_2_2(or_1770_cse, or_1812_nl, fsm_output(3));
  nor_979_nl <= NOT((fsm_output(6)) OR mux_855_nl);
  and_1564_nl <= (fsm_output(6)) AND (fsm_output(3)) AND (fsm_output(5)) AND (NOT
      or_tmp_757);
  mux_856_ssc <= MUX_s_1_2_2(nor_979_nl, and_1564_nl, fsm_output(7));
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_or_1_cse <= and_dcpl_257 OR and_dcpl_265;
  mux_859_nl <= MUX_s_1_2_2(mux_tmp_87, and_1771_cse, fsm_output(1));
  mux_860_nl <= MUX_s_1_2_2(mux_859_nl, nor_tmp_289, fsm_output(0));
  mux_861_nl <= MUX_s_1_2_2(mux_860_nl, (fsm_output(4)), fsm_output(3));
  and_339_ssc <= (NOT mux_861_nl) AND and_dcpl_298;
  mux_863_nl <= MUX_s_1_2_2((NOT nor_tmp_291), nor_tmp_282, fsm_output(5));
  mux_864_nl <= MUX_s_1_2_2(mux_863_nl, mux_tmp_91, fsm_output(3));
  and_343_itm <= (NOT mux_864_nl) AND and_dcpl_308;
  rms_norm_16_div_cmp_b <= reg_rms_norm_16_div_cmp_b_ftd_59_38 & reg_rms_norm_16_div_cmp_b_ftd_37_0
      & reg_rms_norm_16_div_cmp_b_ftd_1;
  rms_norm_16_div_cmp_a <= reg_rms_norm_16_div_cmp_a_ftd & reg_rms_norm_16_div_cmp_a_ftd_1_15_8
      & reg_rms_norm_16_div_cmp_a_ftd_1_7 & reg_rms_norm_16_div_cmp_a_ftd_1_6 & reg_rms_norm_16_div_cmp_a_ftd_1_5
      & reg_rms_norm_16_div_cmp_a_ftd_1_4 & reg_rms_norm_16_div_cmp_a_ftd_1_3 & reg_rms_norm_16_div_cmp_a_ftd_1_2
      & reg_rms_norm_16_div_cmp_a_ftd_1_1 & reg_rms_norm_16_div_cmp_a_ftd_1_0 & STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000");
  and_362_ssc <= and_dcpl_322 AND and_dcpl_319 AND reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      AND (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  nor_907_nl <= NOT((fsm_output(3)) OR (fsm_output(5)) OR (fsm_output(0)) OR (fsm_output(1))
      OR (fsm_output(2)) OR (fsm_output(4)) OR (NOT (fsm_output(8))));
  mux_873_nl <= MUX_s_1_2_2((fsm_output(8)), nor_907_nl, fsm_output(6));
  mux_870_nl <= MUX_s_1_2_2(or_tmp_757, (fsm_output(8)), fsm_output(5));
  or_85_nl <= nor_646_cse OR (fsm_output(8));
  mux_871_nl <= MUX_s_1_2_2(mux_870_nl, or_85_nl, fsm_output(3));
  mux_872_nl <= MUX_s_1_2_2(mux_871_nl, (fsm_output(8)), fsm_output(6));
  mux_874_nl <= MUX_s_1_2_2((NOT mux_873_nl), mux_872_nl, fsm_output(7));
  apply_rotary_pos_emb_1_4_4_rotated_q_and_3_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND mux_874_nl;
  nor_294_nl <= NOT((NOT (fsm_output(4))) OR reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      OR reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      OR (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1));
  mux_876_nl <= MUX_s_1_2_2(nor_tmp_117, mux_tmp_363, nor_294_nl);
  mux_877_nl <= MUX_s_1_2_2(and_1455_cse, mux_876_nl, fsm_output(0));
  mux_878_nl <= MUX_s_1_2_2(mux_877_nl, nor_tmp_117, or_1835_cse);
  apply_rotary_pos_emb_1_4_4_rotated_k_and_6_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND mux_878_nl;
  or_1840_nl <= (NOT (fsm_output(4))) OR reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      OR reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 OR (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd)
      OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  mux_880_nl <= MUX_s_1_2_2(mux_tmp_363, nor_tmp_117, or_1840_nl);
  mux_881_nl <= MUX_s_1_2_2(and_1455_cse, mux_880_nl, fsm_output(0));
  mux_882_nl <= MUX_s_1_2_2(mux_881_nl, nor_tmp_117, or_1835_cse);
  apply_rotary_pos_emb_1_4_4_rotated_k_and_7_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND mux_882_nl;
  nor_301_nl <= NOT((NOT (fsm_output(4))) OR reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      OR reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 OR (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd)
      OR (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1));
  mux_884_nl <= MUX_s_1_2_2(nor_tmp_117, mux_tmp_363, nor_301_nl);
  mux_885_nl <= MUX_s_1_2_2(and_1455_cse, mux_884_nl, fsm_output(0));
  mux_886_nl <= MUX_s_1_2_2(mux_885_nl, nor_tmp_117, or_1835_cse);
  apply_rotary_pos_emb_1_4_4_rotated_k_and_8_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND mux_886_nl;
  or_1848_cse <= (NOT (fsm_output(1))) OR (NOT (fsm_output(0))) OR (fsm_output(8));
  or_1851_cse <= (fsm_output(5)) OR (fsm_output(8));
  nor_305_cse <= NOT((fsm_output(5)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(0))));
  ATTN_2D_LOOP_3_mux_16_itm <= MUX_s_1_16_2((apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2(39)),
      (attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2(39)), (attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2(39)),
      attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_39, (attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2(39)),
      (attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2(39)), (attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2(39)),
      (attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2(39)), (attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2(39)),
      (attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2(39)), (attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2(39)),
      (attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2(39)), (attention_2_1_16_16_4_4_attn_output_3_0_0_sva_2(39)),
      (attention_2_1_16_16_4_4_attn_output_3_0_1_sva_2(39)), (attention_2_1_16_16_4_4_attn_output_3_0_2_sva_2(39)),
      (attention_2_1_16_16_4_4_attn_output_3_0_3_sva_2(39)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  ATTN_2D_LOOP_3_mux_17_itm <= MUX_v_39_16_2((apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2(38
      DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2(38 DOWNTO 0)),
      (attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2(38 DOWNTO 0)), attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_38_0,
      (attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2(38 DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2(38
      DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2(38 DOWNTO 0)),
      (attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2(38 DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2(38
      DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2(38 DOWNTO 0)),
      (attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2(38 DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2(38
      DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_3_0_0_sva_2(38 DOWNTO 0)),
      (attention_2_1_16_16_4_4_attn_output_3_0_1_sva_2(38 DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_3_0_2_sva_2(38
      DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_3_0_3_sva_2(38 DOWNTO 0)),
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  or_1880_cse <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 OR reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  and_28_cse <= (input_0_0_sva_2(39)) AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  or_1879_cse <= (fsm_output(4)) OR (fsm_output(6));
  or_1867_cse <= (NOT (fsm_output(1))) OR (fsm_output(4));
  GEMM_3D_FLOAT_LOOP_4_1_mux1h_5_itm <= MUX_v_40_12_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_1, attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_1,
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_1, attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_1,
      attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_1, attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_1,
      attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_1, attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_1,
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_1, attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_1,
      attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_1, STD_LOGIC_VECTOR'( reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2));
  or_3156_nl <= (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(1)));
  or_3157_nl <= (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (fsm_output(1));
  mux_905_nl <= MUX_s_1_2_2(or_3156_nl, or_3157_nl, fsm_output(7));
  and_404_itm <= (NOT(mux_905_nl OR (fsm_output(8)))) AND and_dcpl_364 AND and_dcpl_194;
  rms_norm_16_variance_or_1_cse <= and_dcpl_242 OR (and_dcpl_239 AND and_dcpl_182);
  nor_985_nl <= NOT((fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(5)) OR (fsm_output(0))
      OR (fsm_output(1)) OR (fsm_output(2)));
  and_1566_nl <= (fsm_output(3)) AND (fsm_output(5)) AND (fsm_output(0)) AND (fsm_output(1))
      AND (NOT (fsm_output(2)));
  nor_986_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(5)) OR (fsm_output(0)) OR
      (fsm_output(1)) OR (NOT (fsm_output(2))));
  mux_947_nl <= MUX_s_1_2_2(and_1566_nl, nor_986_nl, fsm_output(6));
  mux_948_nl <= MUX_s_1_2_2(nor_985_nl, mux_947_nl, fsm_output(7));
  GEMM_3D_FLOAT_LOOP_4_1_nand_itm <= NOT(mux_948_nl AND and_dcpl_61);
  mux_941_nl <= MUX_s_1_2_2(mux_tmp_916, or_1197_cse, fsm_output(4));
  mux_939_nl <= MUX_s_1_2_2(mux_tmp_936, or_1197_cse, fsm_output(4));
  mux_940_nl <= MUX_s_1_2_2(mux_939_nl, mux_tmp_937, or_1880_cse);
  mux_942_nl <= MUX_s_1_2_2(mux_941_nl, mux_940_nl, fsm_output(0));
  mux_938_nl <= MUX_s_1_2_2(mux_tmp_937, mux_tmp_922, fsm_output(0));
  mux_943_nl <= MUX_s_1_2_2(mux_942_nl, mux_938_nl, fsm_output(1));
  mux_933_nl <= MUX_s_1_2_2(or_tmp_808, or_tmp_805, fsm_output(4));
  mux_934_nl <= MUX_s_1_2_2(mux_933_nl, mux_tmp_927, fsm_output(0));
  mux_932_nl <= MUX_s_1_2_2(or_tmp_805, or_tmp_812, fsm_output(4));
  mux_935_nl <= MUX_s_1_2_2(mux_934_nl, mux_932_nl, fsm_output(1));
  mux_944_nl <= MUX_s_1_2_2(mux_943_nl, mux_935_nl, fsm_output(5));
  mux_928_nl <= MUX_s_1_2_2(or_362_cse, or_361_cse, or_1879_cse);
  mux_929_nl <= MUX_s_1_2_2(mux_928_nl, mux_tmp_927, fsm_output(0));
  mux_930_nl <= MUX_s_1_2_2(mux_tmp_915, mux_929_nl, fsm_output(1));
  mux_931_nl <= MUX_s_1_2_2(mux_tmp_908, mux_930_nl, fsm_output(5));
  mux_945_nl <= MUX_s_1_2_2(mux_944_nl, mux_931_nl, fsm_output(3));
  mux_920_nl <= MUX_s_1_2_2(mux_tmp_919, or_tmp_813, fsm_output(4));
  mux_923_nl <= MUX_s_1_2_2(mux_tmp_922, mux_920_nl, fsm_output(0));
  mux_917_nl <= MUX_s_1_2_2(mux_tmp_916, or_tmp_813, fsm_output(4));
  mux_918_nl <= MUX_s_1_2_2(mux_917_nl, mux_tmp_910, fsm_output(0));
  mux_924_nl <= MUX_s_1_2_2(mux_923_nl, mux_918_nl, fsm_output(1));
  mux_925_nl <= MUX_s_1_2_2(mux_924_nl, mux_tmp_915, fsm_output(5));
  mux_912_nl <= MUX_s_1_2_2(mux_tmp_908, mux_tmp_910, fsm_output(0));
  mux_911_nl <= MUX_s_1_2_2(mux_tmp_910, mux_tmp_908, fsm_output(0));
  mux_913_nl <= MUX_s_1_2_2(mux_912_nl, mux_911_nl, fsm_output(1));
  mux_907_nl <= MUX_s_1_2_2(mux_tmp_906, or_tmp_805, or_1867_cse);
  mux_914_nl <= MUX_s_1_2_2(mux_913_nl, mux_907_nl, fsm_output(5));
  mux_926_nl <= MUX_s_1_2_2(mux_925_nl, mux_914_nl, fsm_output(3));
  mux_946_nl <= MUX_s_1_2_2(mux_945_nl, mux_926_nl, fsm_output(2));
  GEMM_3D_FLOAT_LOOP_4_1_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND mux_946_nl;
  or_1907_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01"));
  and_1572_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"));
  or_1908_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"));
  and_1570_cse <= (fsm_output(1)) AND (fsm_output(2)) AND (fsm_output(4));
  nor_992_cse <= NOT((fsm_output(2)) OR (fsm_output(4)));
  nand_240_cse <= NOT((fsm_output(1)) AND (fsm_output(0)) AND (fsm_output(2)) AND
      (fsm_output(4)));
  mux_958_cse <= MUX_s_1_2_2(or_tmp_48, or_133_cse, fsm_output(5));
  or_1890_nl <= (fsm_output(3)) OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR (fsm_output(6));
  or_3158_nl <= (NOT (fsm_output(2))) OR (fsm_output(6));
  nand_318_nl <= NOT((fsm_output(2)) AND (fsm_output(6)));
  mux_950_nl <= MUX_s_1_2_2(or_3158_nl, nand_318_nl, fsm_output(0));
  or_1889_nl <= (NOT (fsm_output(3))) OR (fsm_output(5)) OR mux_950_nl;
  mux_951_nl <= MUX_s_1_2_2(or_1890_nl, or_1889_nl, fsm_output(7));
  nor_990_nl <= NOT((fsm_output(8)) OR mux_951_nl);
  nor_988_nl <= NOT(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4 OR (NOT (fsm_output(0)))
      OR (fsm_output(2)) OR (fsm_output(6)));
  nor_989_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(6)));
  mux_949_nl <= MUX_s_1_2_2(nor_988_nl, nor_989_nl, fsm_output(5));
  and_1568_nl <= (NOT((NOT (fsm_output(8))) OR (fsm_output(7)) OR (NOT (fsm_output(3)))))
      AND mux_949_nl;
  mux_952_nl <= MUX_s_1_2_2(nor_990_nl, and_1568_nl, fsm_output(4));
  and_416_itm <= mux_952_nl AND (fsm_output(1));
  nand_47_nl <= NOT((fsm_output(5)) AND nor_998_cse);
  mux_985_nl <= MUX_s_1_2_2(nand_47_nl, or_tmp_798, fsm_output(3));
  and_428_itm <= (NOT mux_985_nl) AND and_dcpl_390;
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_cse <= and_dcpl_382 OR and_dcpl_386;
  or_3206_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("110"));
  or_3207_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("001"));
  mux_2236_nl <= MUX_s_1_2_2(or_3206_nl, or_3207_nl, fsm_output(6));
  nor_1314_cse <= NOT(mux_2236_nl OR (fsm_output(8)));
  or_1923_nl <= (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(8));
  or_1922_nl <= (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(8)));
  mux_978_nl <= MUX_s_1_2_2(or_1923_nl, or_1922_nl, fsm_output(4));
  or_1920_nl <= (fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(8));
  mux_979_nl <= MUX_s_1_2_2(mux_978_nl, or_1920_nl, fsm_output(2));
  or_1919_nl <= (NOT (fsm_output(4))) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR (fsm_output(8));
  or_1918_nl <= (fsm_output(4)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(8));
  mux_977_nl <= MUX_s_1_2_2(or_1919_nl, or_1918_nl, fsm_output(2));
  mux_980_nl <= MUX_s_1_2_2(mux_979_nl, mux_977_nl, fsm_output(7));
  or_3159_nl <= (fsm_output(1)) OR mux_980_nl;
  or_1916_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(8));
  nand_321_nl <= NOT(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4 AND (fsm_output(3))
      AND (NOT (fsm_output(6))) AND (fsm_output(8)));
  mux_976_nl <= MUX_s_1_2_2(or_1916_nl, nand_321_nl, fsm_output(4));
  or_3160_nl <= (NOT (fsm_output(1))) OR (fsm_output(7)) OR (fsm_output(2)) OR mux_976_nl;
  mux_981_nl <= MUX_s_1_2_2(or_3159_nl, or_3160_nl, fsm_output(0));
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_5_itm <= mux_981_nl OR (fsm_output(5));
  mux_969_nl <= MUX_s_1_2_2(or_tmp_48, or_133_cse, and_1559_cse);
  mux_970_nl <= MUX_s_1_2_2(mux_969_nl, mux_tmp_968, fsm_output(0));
  nor_991_nl <= NOT(and_1570_cse OR (fsm_output(8)));
  mux_971_nl <= MUX_s_1_2_2(mux_970_nl, nor_991_nl, fsm_output(5));
  mux_964_nl <= MUX_s_1_2_2(and_dcpl_61, mux_528_cse, or_1908_cse);
  mux_963_nl <= MUX_s_1_2_2(and_dcpl_61, mux_528_cse, or_1907_cse);
  mux_965_nl <= MUX_s_1_2_2(mux_964_nl, mux_963_nl, fsm_output(0));
  nand_319_nl <= NOT((NOT((fsm_output(1)) AND (fsm_output(2)) AND (fsm_output(4))))
      AND (fsm_output(8)));
  mux_961_nl <= MUX_s_1_2_2(mux_tmp_960, nand_319_nl, fsm_output(0));
  mux_966_nl <= MUX_s_1_2_2((NOT mux_965_nl), mux_961_nl, fsm_output(5));
  mux_972_nl <= MUX_s_1_2_2(mux_971_nl, mux_966_nl, fsm_output(3));
  or_1901_nl <= nor_992_cse OR (fsm_output(8));
  or_1899_nl <= and_1572_cse OR (fsm_output(4)) OR (fsm_output(8));
  mux_957_nl <= MUX_s_1_2_2(or_1901_nl, or_1899_nl, fsm_output(5));
  mux_959_nl <= MUX_s_1_2_2(mux_958_cse, mux_957_nl, fsm_output(3));
  mux_973_nl <= MUX_s_1_2_2(mux_972_nl, mux_959_nl, fsm_output(6));
  or_1898_nl <= (fsm_output(2)) OR (fsm_output(4)) OR (fsm_output(8));
  mux_954_nl <= MUX_s_1_2_2(or_1898_nl, or_tmp_833, or_1732_cse);
  mux_955_nl <= MUX_s_1_2_2(or_tmp_757, mux_954_nl, fsm_output(5));
  or_1895_nl <= (fsm_output(5)) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_956_nl <= MUX_s_1_2_2(mux_955_nl, or_1895_nl, fsm_output(3));
  nand_46_nl <= NOT((fsm_output(6)) AND (NOT mux_956_nl));
  mux_974_nl <= MUX_s_1_2_2(mux_973_nl, nand_46_nl, fsm_output(7));
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND mux_974_nl;
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_7_cse <= and_dcpl_328 AND and_428_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_8_cse <= and_dcpl_313 AND and_428_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_9_cse <= and_dcpl_587 AND and_dcpl_190 AND
      and_428_itm;
  compute_sqrt_for_i_and_2_cse <= (NOT and_dcpl_557) AND and_dcpl_414;
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c0 OR and_dcpl_242 OR
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c2 OR LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c3
      OR LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c5 OR and_dcpl_410 OR LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c7
      OR and_dcpl_414);
  compute_sqrt_for_i_and_cse <= and_dcpl_201 AND and_1474_cse AND and_dcpl_199 AND
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c7;
  nor_1311_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR or_dcpl_1050);
  mux_2227_nl <= MUX_s_1_2_2(nor_1311_nl, mux_tmp_1451, fsm_output(5));
  mux_2228_nl <= MUX_s_1_2_2(mux_2227_nl, and_tmp_42, fsm_output(3));
  mux_2229_nl <= MUX_s_1_2_2(mux_2228_nl, (NOT or_tmp_755), fsm_output(6));
  compute_sqrt_for_i_and_4_cse <= mux_2229_nl AND and_dcpl_295 AND LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c7;
  compute_sqrt_for_i_and_5_cse <= (and_dcpl_328 OR and_dcpl_635) AND LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c7;
  and_1773_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"));
  or_1983_cse <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  or_1985_cse <= CONV_SL_1_1(fsm_output(7 DOWNTO 5)/=STD_LOGIC_VECTOR'("011"));
  or_1984_cse <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  nor_1026_cse <= NOT((fsm_output(0)) OR (fsm_output(5)));
  for_for_and_13_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (and_dcpl_415
      OR for_for_strm_in_tmp_sva_31_2_mx0c1);
  and_474_rgt <= and_dcpl_342 AND and_dcpl_336 AND and_dcpl_433;
  and_476_rgt <= or_dcpl_1071 AND and_dcpl_185 AND and_dcpl_422;
  and_480_rgt <= and_dcpl_350 AND and_dcpl_190;
  for_for_and_14_rgt <= (NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd OR reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1))
      AND and_dcpl_442;
  for_for_and_15_rgt <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd)
      AND and_dcpl_442;
  for_for_and_16_rgt <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1)
      AND and_dcpl_442;
  for_for_and_17_rgt <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      AND and_dcpl_442;
  and_485_rgt <= and_dcpl_241 AND (fsm_output(5)) AND SOFTMAX_LOOP_3_acc_3_itm_40_1
      AND (fsm_output(3)) AND and_dcpl_45;
  and_486_rgt <= and_dcpl_376 AND and_dcpl_221;
  for_for_or_1_rgt <= and_dcpl_448 OR (and_dcpl_449 AND and_dcpl_200 AND and_dcpl_261);
  nand_328_nl <= NOT((fsm_output(2)) AND (fsm_output(5)) AND (fsm_output(3)) AND
      (fsm_output(7)));
  or_2016_nl <= (fsm_output(5)) OR (fsm_output(3)) OR (fsm_output(7));
  or_2015_nl <= SOFTMAX_LOOP_3_acc_3_itm_40_1 OR not_tmp_549;
  mux_1068_nl <= MUX_s_1_2_2(or_2016_nl, or_2015_nl, fsm_output(0));
  or_2014_nl <= (fsm_output(0)) OR not_tmp_549;
  mux_1069_nl <= MUX_s_1_2_2(mux_1068_nl, or_2014_nl, fsm_output(2));
  mux_1070_nl <= MUX_s_1_2_2(nand_328_nl, mux_1069_nl, fsm_output(1));
  or_2013_nl <= (NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 OR reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1))
      OR (NOT (fsm_output(0))) OR (fsm_output(5)) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1066_nl <= MUX_s_1_2_2(or_2013_nl, or_tmp_938, fsm_output(2));
  or_2007_nl <= (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_2006_nl <= (fsm_output(3)) OR (fsm_output(7));
  mux_1064_nl <= MUX_s_1_2_2(or_2007_nl, or_2006_nl, fsm_output(5));
  or_2008_nl <= (fsm_output(0)) OR mux_1064_nl;
  mux_1065_nl <= MUX_s_1_2_2(or_tmp_938, or_2008_nl, fsm_output(2));
  mux_1067_nl <= MUX_s_1_2_2(mux_1066_nl, mux_1065_nl, fsm_output(1));
  mux_1071_nl <= MUX_s_1_2_2(mux_1070_nl, mux_1067_nl, fsm_output(4));
  nand_329_nl <= NOT((fsm_output(4)) AND (NOT (fsm_output(1))) AND (fsm_output(2))
      AND (fsm_output(0)) AND (fsm_output(5)) AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_1072_nl <= MUX_s_1_2_2(mux_1071_nl, nand_329_nl, fsm_output(6));
  QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (mux_1072_nl OR (fsm_output(8)));
  and_37_cse <= (RMS_NORM_LOOP_2_2_i_4_0_sva_1(4)) AND reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_8_seb <= NOT(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva_mx0w3
      AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  mux_1114_nl <= MUX_s_1_2_2((NOT nor_tmp_289), mux_tmp_1113, fsm_output(0));
  mux_1115_nl <= MUX_s_1_2_2(mux_1114_nl, or_tmp_992, fsm_output(6));
  mux_1116_nl <= MUX_s_1_2_2(or_tmp_993, mux_1115_nl, fsm_output(7));
  apply_rotary_pos_emb_1_4_4_rotated_q_and_37_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT or_dcpl_1068) OR apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c0
      OR apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c1 OR and_dcpl_477 OR
      and_dcpl_220 OR and_dcpl_222 OR and_dcpl_187) AND (NOT((NOT mux_1116_nl) AND
      and_dcpl_478));
  or_2081_nl <= (fsm_output(1)) OR or_dcpl_1050;
  or_2080_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (NOT (fsm_output(4)));
  mux_1117_nl <= MUX_s_1_2_2(or_2081_nl, or_2080_nl, fsm_output(0));
  mux_1118_nl <= MUX_s_1_2_2(mux_1117_nl, or_tmp_992, fsm_output(6));
  mux_1119_nl <= MUX_s_1_2_2(or_tmp_993, mux_1118_nl, fsm_output(7));
  attention_2_1_16_16_4_4_attn_output_and_25_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT((NOT mux_1119_nl) AND and_dcpl_478));
  or_3212_tmp <= (and_dcpl_1233 AND GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva_mx0w0)
      OR mux_tmp_1163;
  or_3213_tmp <= (and_dcpl_1233 AND GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva_mx0w0)
      OR mux_tmp_1163;
  or_3214_tmp <= (and_dcpl_1233 AND GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva_mx0w0)
      OR attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c10;
  nor_366_cse <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")));
  or_3167_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("10"));
  or_2154_cse <= (NOT (fsm_output(5))) OR (fsm_output(7));
  nor_1044_cse <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(2)))
      OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1045_cse <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(1))
      OR (NOT (fsm_output(2))) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1208_nl <= MUX_s_1_2_2(and_dcpl_449, and_dcpl_263, fsm_output(1));
  mux_1209_nl <= MUX_s_1_2_2(and_dcpl_341, mux_1208_nl, fsm_output(3));
  mux_1210_nl <= MUX_s_1_2_2(mux_1209_nl, nor_1044_cse, fsm_output(6));
  mux_1211_nl <= MUX_s_1_2_2(mux_1210_nl, nor_1045_cse, fsm_output(7));
  and_581_ssc <= mux_1211_nl AND and_dcpl_338;
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_nand_seb <= NOT(and_dcpl_381 AND nor_777_cse AND
      and_dcpl_198);
  nor_1046_nl <= NOT((fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(1)) OR (NOT
      (fsm_output(2))));
  and_1597_nl <= (fsm_output(6)) AND (fsm_output(0)) AND (fsm_output(1)) AND (NOT
      (fsm_output(2)));
  mux_1212_nl <= MUX_s_1_2_2(nor_1046_nl, and_1597_nl, fsm_output(7));
  and_585_seb <= mux_1212_nl AND and_dcpl_201 AND and_dcpl_189;
  mux_1231_nl <= MUX_s_1_2_2(mux_tmp_1229, mux_tmp_1219, fsm_output(1));
  mux_1230_nl <= MUX_s_1_2_2(mux_tmp_1229, mux_tmp_1219, fsm_output(2));
  mux_1232_nl <= MUX_s_1_2_2(mux_1231_nl, mux_1230_nl, fsm_output(0));
  mux_1233_nl <= MUX_s_1_2_2(mux_1232_nl, or_1795_cse, fsm_output(6));
  mux_1226_nl <= MUX_s_1_2_2(mux_tmp_1218, or_tmp_1051, fsm_output(2));
  mux_1225_nl <= MUX_s_1_2_2(mux_tmp_1218, or_2154_cse, fsm_output(2));
  mux_1227_nl <= MUX_s_1_2_2(mux_1226_nl, mux_1225_nl, or_1732_cse);
  or_2152_nl <= (NOT((fsm_output(2)) OR (NOT (fsm_output(7))))) OR (fsm_output(8));
  or_2151_nl <= (NOT((fsm_output(2)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7)))))
      OR (fsm_output(8));
  mux_1223_nl <= MUX_s_1_2_2(or_2152_nl, or_2151_nl, fsm_output(1));
  or_2150_nl <= (or_3167_cse AND (fsm_output(5)) AND (fsm_output(7))) OR (fsm_output(8));
  mux_1224_nl <= MUX_s_1_2_2(mux_1223_nl, or_2150_nl, fsm_output(0));
  mux_1228_nl <= MUX_s_1_2_2(mux_1227_nl, mux_1224_nl, fsm_output(6));
  mux_1234_nl <= MUX_s_1_2_2(mux_1233_nl, mux_1228_nl, fsm_output(4));
  mux_1220_nl <= MUX_s_1_2_2(mux_tmp_1219, mux_tmp_1218, and_1559_cse);
  or_2145_nl <= (NOT (fsm_output(2))) OR (fsm_output(5));
  mux_1216_nl <= MUX_s_1_2_2(or_361_cse, or_362_cse, or_2145_nl);
  mux_1217_nl <= MUX_s_1_2_2(or_1795_cse, mux_1216_nl, nor_366_cse);
  mux_1221_nl <= MUX_s_1_2_2(mux_1220_nl, mux_1217_nl, fsm_output(6));
  or_2142_nl <= (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(8)));
  mux_1213_nl <= MUX_s_1_2_2(or_tmp_1051, or_2142_nl, fsm_output(1));
  or_2140_nl <= and_1559_cse OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT
      (fsm_output(8)));
  mux_1214_nl <= MUX_s_1_2_2(mux_1213_nl, or_2140_nl, fsm_output(0));
  or_2138_nl <= ((fsm_output(5)) AND (fsm_output(7))) OR (fsm_output(8));
  mux_1215_nl <= MUX_s_1_2_2(mux_1214_nl, or_2138_nl, fsm_output(6));
  mux_1222_nl <= MUX_s_1_2_2(mux_1221_nl, mux_1215_nl, fsm_output(4));
  mux_1235_nl <= MUX_s_1_2_2(mux_1234_nl, mux_1222_nl, fsm_output(3));
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_1_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND mux_1235_nl;
  attention_abs_qelse_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT(((and_1637_cse OR (fsm_output(3))) XOR (fsm_output(4))) AND and_dcpl_270));
  compute_sqrt_guess_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((and_dcpl_192 AND and_dcpl_209) OR and_dcpl_290);
  nor_1229_cse <= NOT(reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  and_1191_rgt <= and_dcpl_1061 AND and_dcpl_45 AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      AND nor_1229_cse AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd;
  mux_1310_nl <= MUX_s_1_2_2(or_tmp_611, or_tmp_1128, fsm_output(3));
  and_622_rgt <= (NOT mux_1310_nl) AND and_dcpl_581;
  operator_40_24_true_AC_TRN_AC_WRAP_1_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT(or_dcpl_1040 AND and_dcpl_191 AND and_dcpl_321 AND and_dcpl_1141));
  operator_40_24_true_AC_TRN_AC_WRAP_1_conc_1_itm_11_0 <= MUX_v_12_16_2(STD_LOGIC_VECTOR'(
      "011110001010"), STD_LOGIC_VECTOR'( "011101010010"), STD_LOGIC_VECTOR'( "100000010100"),
      STD_LOGIC_VECTOR'( "011100010010"), STD_LOGIC_VECTOR'( "011100110010"), STD_LOGIC_VECTOR'(
      "100000011110"), STD_LOGIC_VECTOR'( "011101100011"), STD_LOGIC_VECTOR'( "100000101100"),
      STD_LOGIC_VECTOR'( "011111110100"), STD_LOGIC_VECTOR'( "011100010000"), STD_LOGIC_VECTOR'(
      "011110000101"), STD_LOGIC_VECTOR'( "100001110110"), STD_LOGIC_VECTOR'( "011101111110"),
      STD_LOGIC_VECTOR'( "011110001010"), STD_LOGIC_VECTOR'( "100000111010"), STD_LOGIC_VECTOR'(
      "100001001110"), reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  operator_40_24_true_AC_TRN_AC_WRAP_1_conc_3_itm_8_0 <= MUX_v_9_16_2(STD_LOGIC_VECTOR'(
      "011001100"), STD_LOGIC_VECTOR'( "001101100"), STD_LOGIC_VECTOR'( "101011100"),
      STD_LOGIC_VECTOR'( "100110000"), STD_LOGIC_VECTOR'( "010100011"), STD_LOGIC_VECTOR'(
      "101100000"), STD_LOGIC_VECTOR'( "011001100"), STD_LOGIC_VECTOR'( "101000111"),
      STD_LOGIC_VECTOR'( "110000011"), STD_LOGIC_VECTOR'( "010111100"), STD_LOGIC_VECTOR'(
      "010001100"), STD_LOGIC_VECTOR'( "100000000"), STD_LOGIC_VECTOR'( "011000000"),
      STD_LOGIC_VECTOR'( "000100111"), STD_LOGIC_VECTOR'( "110111000"), STD_LOGIC_VECTOR'(
      "101110011"), reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  or_3174_nl <= (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  nand_344_nl <= NOT((fsm_output(6)) AND (fsm_output(3)) AND (fsm_output(2)));
  mux_1308_nl <= MUX_s_1_2_2(or_3174_nl, nand_344_nl, fsm_output(7));
  and_615_itm <= (NOT(mux_1308_nl OR (fsm_output(8)))) AND and_1651_cse AND nor_1026_cse;
  operator_40_24_true_AC_TRN_AC_WRAP_1_and_4_cse <= (NOT and_1191_rgt) AND and_622_rgt;
  attention_2_1_16_16_4_4_quantized_hidden_states_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1087 OR and_dcpl_618)) OR or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_cse <= QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1
      AND and_dcpl_619;
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_cse <= (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1)
      AND and_dcpl_619;
  attention_2_1_16_16_4_4_quantized_hidden_states_and_1_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1086 OR and_dcpl_618)) OR or_dcpl_1104);
  attention_2_1_16_16_4_4_quantized_hidden_states_and_2_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1067 OR and_dcpl_618)) OR or_dcpl_1104);
  attention_2_1_16_16_4_4_quantized_hidden_states_and_3_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1079 OR and_dcpl_618)) OR or_dcpl_1104);
  or_3185_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  and_1637_cse <= or_1732_cse AND (fsm_output(2));
  RMS_NORM_LOOP_2_2_i_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (and_dcpl_477 OR RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c1 OR and_dcpl_410
      OR and_dcpl_620 OR RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c4 OR and_dcpl_255);
  RMS_NORM_LOOP_2_2_i_and_9_cse <= and_dcpl_564 AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1)
      AND and_dcpl_620;
  or_2249_cse <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  and_633_itm <= and_dcpl_588 AND and_dcpl_592;
  and_654_itm <= and_dcpl_588 AND and_dcpl_613;
  and_648_itm <= and_dcpl_588 AND and_dcpl_607;
  and_642_itm <= and_dcpl_588 AND and_dcpl_601;
  and_636_itm <= and_dcpl_588 AND and_dcpl_595;
  and_629_itm <= and_dcpl_588 AND and_dcpl_586;
  and_639_itm <= and_dcpl_588 AND and_dcpl_598;
  and_645_itm <= and_dcpl_588 AND and_dcpl_604;
  and_651_itm <= and_dcpl_588 AND and_dcpl_610;
  and_657_itm <= and_dcpl_588 AND and_dcpl_616;
  and_1638_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111"));
  nor_1106_cse <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
  and_937_ssc <= (NOT(mux_tmp_1426 OR (fsm_output(8)))) AND and_dcpl_338 AND and_dcpl_45;
  nand_71_nl <= NOT((fsm_output(6)) AND (fsm_output(3)) AND (NOT(and_1474_cse OR
      (NOT (fsm_output(2))) OR (fsm_output(4)))));
  mux_1636_nl <= MUX_s_1_2_2(or_tmp_1221, or_tmp_1128, fsm_output(0));
  mux_1637_nl <= MUX_s_1_2_2(or_tmp_1203, mux_1636_nl, fsm_output(3));
  or_2563_nl <= (fsm_output(6)) OR mux_1637_nl;
  mux_1638_nl <= MUX_s_1_2_2(nand_71_nl, or_2563_nl, fsm_output(7));
  nor_1324_seb <= NOT(mux_1638_nl OR or_1851_cse);
  and_679_nl <= (fsm_output(5)) AND mux_tmp_1451;
  mux_1452_nl <= MUX_s_1_2_2(and_679_nl, and_tmp_42, fsm_output(3));
  mux_1453_nl <= MUX_s_1_2_2(mux_1452_nl, (NOT or_tmp_755), fsm_output(6));
  CACHE_UPDATE_LOOP_3_k_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT(mux_1453_nl AND and_dcpl_295));
  QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_or_cse <= and_dcpl_888
      OR (and_dcpl_362 AND and_dcpl_237);
  nand_197_cse <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")));
  nor_777_cse <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  nand_350_nl <= NOT(or_2500_cse AND (fsm_output(7)));
  or_2355_nl <= (fsm_output(1)) OR (NOT (fsm_output(7)));
  mux_1456_nl <= MUX_s_1_2_2(nand_350_nl, or_2355_nl, fsm_output(0));
  nor_1115_nl <= NOT((fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR mux_1456_nl);
  nor_1116_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(0))
      OR (fsm_output(1)) OR (fsm_output(7)));
  nor_1114_nl <= NOT(nor_777_cse OR (fsm_output(7)));
  mux_1454_nl <= MUX_s_1_2_2(nor_1114_nl, (fsm_output(7)), fsm_output(6));
  nor_1117_nl <= NOT((fsm_output(3)) OR (NOT mux_1454_nl));
  mux_1455_nl <= MUX_s_1_2_2(nor_1116_nl, nor_1117_nl, fsm_output(2));
  mux_1457_nl <= MUX_s_1_2_2(nor_1115_nl, mux_1455_nl, fsm_output(5));
  GEMM_3D_FLOAT_LOOP_1_i_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((mux_1457_nl AND and_dcpl_201) OR GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c1
      OR GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c2);
  nand_126_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 3)=STD_LOGIC_VECTOR'("111")));
  mux_1490_nl <= MUX_s_1_2_2(nand_126_nl, mux_tmp_1489, fsm_output(6));
  input_and_28_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT((NOT
      mux_1490_nl) AND and_dcpl_26));
  and_699_ssc <= or_dcpl_1116 AND and_dcpl_202 AND and_dcpl_642;
  and_745_ssc <= or_dcpl_1131 AND and_dcpl_202 AND and_dcpl_642;
  or_2456_cse <= (fsm_output(6)) OR (NOT (fsm_output(8)));
  or_2457_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001"));
  or_2455_cse <= (fsm_output(6)) OR (fsm_output(8));
  or_2460_cse <= (fsm_output(4)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(6)))
      OR (fsm_output(8));
  or_2451_cse <= (fsm_output(4)) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (fsm_output(8));
  mux_1522_cse <= MUX_s_1_2_2(or_2456_cse, or_2455_cse, fsm_output(7));
  or_2443_nl <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (fsm_output(4));
  mux_1513_cse <= MUX_s_1_2_2(or_2443_nl, or_tmp_1128, fsm_output(0));
  mux_1496_nl <= MUX_s_1_2_2(or_tmp_931, or_2154_cse, fsm_output(4));
  or_2429_nl <= (fsm_output(6)) OR mux_1496_nl;
  or_2426_nl <= (fsm_output(2)) OR (NOT (fsm_output(3))) OR (fsm_output(0));
  mux_1497_nl <= MUX_s_1_2_2(or_2429_nl, or_tmp_1291, or_2426_nl);
  nand_354_nl <= NOT((fsm_output(4)) AND (fsm_output(5)) AND (fsm_output(7)));
  mux_1492_nl <= MUX_s_1_2_2(or_tmp_930, nand_354_nl, fsm_output(6));
  mux_1493_nl <= MUX_s_1_2_2(or_tmp_1291, mux_1492_nl, fsm_output(0));
  nand_355_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 4)=STD_LOGIC_VECTOR'("0111")));
  mux_1494_nl <= MUX_s_1_2_2(mux_1493_nl, nand_355_nl, fsm_output(3));
  mux_1495_nl <= MUX_s_1_2_2(or_tmp_1291, mux_1494_nl, fsm_output(2));
  mux_1498_nl <= MUX_s_1_2_2(mux_1497_nl, mux_1495_nl, fsm_output(1));
  nor_1138_m1c <= NOT(mux_1498_nl OR (fsm_output(8)));
  or_2442_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR (NOT
      RESHAPE_2D_TO_3D_LOOP_2_2_and_cse) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(7)))
      OR (fsm_output(6)) OR (fsm_output(8));
  mux_1510_nl <= MUX_s_1_2_2(or_2442_nl, or_tmp_1296, fsm_output(5));
  or_2441_nl <= (NOT RESHAPE_2D_TO_3D_LOOP_2_2_and_cse) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (fsm_output(8));
  mux_1507_nl <= MUX_s_1_2_2(or_2441_nl, mux_tmp_1519, fsm_output(3));
  or_2438_nl <= (NOT (z_out_4(2))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(7)))
      OR (fsm_output(6)) OR (fsm_output(8));
  mux_1505_nl <= MUX_s_1_2_2(or_2438_nl, or_2451_cse, fsm_output(3));
  mux_1508_nl <= MUX_s_1_2_2(mux_1507_nl, mux_1505_nl, fsm_output(2));
  or_2436_nl <= reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("010"));
  mux_1503_nl <= MUX_s_1_2_2(or_2436_nl, or_1197_cse, fsm_output(4));
  mux_1504_nl <= MUX_s_1_2_2(or_2451_cse, mux_1503_nl, fsm_output(3));
  nand_64_nl <= NOT((fsm_output(2)) AND (NOT mux_1504_nl));
  mux_1509_nl <= MUX_s_1_2_2(mux_1508_nl, nand_64_nl, fsm_output(5));
  mux_1511_nl <= MUX_s_1_2_2(mux_1510_nl, mux_1509_nl, fsm_output(1));
  mux_1500_nl <= MUX_s_1_2_2(or_2460_cse, mux_2092_cse, fsm_output(3));
  or_2431_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(7)))
      OR (fsm_output(6)) OR (fsm_output(8));
  mux_1501_nl <= MUX_s_1_2_2(mux_1500_nl, or_2431_nl, fsm_output(2));
  mux_1502_nl <= MUX_s_1_2_2(mux_1501_nl, or_tmp_1296, fsm_output(5));
  nand_63_nl <= NOT((fsm_output(1)) AND (NOT mux_1502_nl));
  mux_1512_itm <= MUX_s_1_2_2(mux_1511_nl, nand_63_nl, fsm_output(0));
  mux_1529_nl <= MUX_s_1_2_2(or_2460_cse, mux_tmp_1519, fsm_output(3));
  or_2459_nl <= (fsm_output(3)) OR mux_tmp_1519;
  mux_1530_nl <= MUX_s_1_2_2(mux_1529_nl, or_2459_nl, fsm_output(0));
  or_2458_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(7))) OR (fsm_output(6))
      OR (fsm_output(8));
  mux_1527_nl <= MUX_s_1_2_2(or_2458_nl, mux_tmp_1519, fsm_output(3));
  mux_1528_nl <= MUX_s_1_2_2(or_tmp_1320, mux_1527_nl, fsm_output(0));
  mux_1531_nl <= MUX_s_1_2_2(mux_1530_nl, mux_1528_nl, fsm_output(1));
  mux_1532_nl <= MUX_s_1_2_2(mux_1531_nl, or_tmp_1316, fsm_output(5));
  mux_1523_nl <= MUX_s_1_2_2(or_2457_cse, mux_1522_cse, fsm_output(4));
  mux_1524_nl <= MUX_s_1_2_2(mux_tmp_1519, mux_1523_nl, fsm_output(3));
  mux_1520_nl <= MUX_s_1_2_2(mux_tmp_1519, or_2451_cse, fsm_output(3));
  mux_1521_nl <= MUX_s_1_2_2(or_tmp_1320, mux_1520_nl, fsm_output(0));
  mux_1525_nl <= MUX_s_1_2_2(mux_1524_nl, mux_1521_nl, fsm_output(1));
  or_2448_nl <= (NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010"));
  mux_1517_nl <= MUX_s_1_2_2(or_tmp_1316, or_2448_nl, fsm_output(0));
  or_2446_nl <= (NOT((NOT((fsm_output(0)) OR (NOT reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1)
      OR (NOT (fsm_output(3))))) OR (fsm_output(4)))) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("010"));
  mux_1518_nl <= MUX_s_1_2_2(mux_1517_nl, or_2446_nl, fsm_output(1));
  mux_1526_nl <= MUX_s_1_2_2(mux_1525_nl, mux_1518_nl, fsm_output(5));
  mux_1533_nl <= MUX_s_1_2_2(mux_1532_nl, mux_1526_nl, fsm_output(2));
  APPLY_ROTARY_POS_EMB_LOOP_1_i_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND mux_1533_nl;
  mux_1540_nl <= MUX_s_1_2_2(not_tmp_699, or_tmp_1132, fsm_output(7));
  mux_1539_nl <= MUX_s_1_2_2(not_tmp_699, or_tmp_1218, fsm_output(7));
  mux_1541_nl <= MUX_s_1_2_2(mux_1540_nl, mux_1539_nl, reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  nor_1144_itm <= NOT(mux_1541_nl OR (fsm_output(8)));
  attention_2_1_16_16_4_4_q_proj_and_4_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((and_dcpl_588 AND and_dcpl_721) OR and_dcpl_240 OR and_dcpl_626);
  attention_2_1_16_16_4_4_v_proj_re_and_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (and_dcpl_619 OR and_dcpl_725 OR and_dcpl_726 OR and_dcpl_410);
  and_1651_cse <= (fsm_output(4)) AND (fsm_output(1));
  or_2480_cse <= (fsm_output(4)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(8));
  mux_1551_cse <= MUX_s_1_2_2(or_tmp_464, or_2456_cse, fsm_output(5));
  or_2481_cse <= and_1651_cse OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(8));
  mux_1559_cse <= MUX_s_1_2_2(nand_tmp_66, mux_tmp_1549, fsm_output(4));
  mux_1557_cse <= MUX_s_1_2_2(mux_tmp_1549, mux_tmp_1548, and_1651_cse);
  and_1652_nl <= (fsm_output(1)) AND (fsm_output(5));
  mux_1554_nl <= MUX_s_1_2_2(mux_tmp_121, or_tmp_464, and_1652_nl);
  mux_1555_cse <= MUX_s_1_2_2(mux_tmp_1549, mux_1554_nl, fsm_output(4));
  mux_1552_nl <= MUX_s_1_2_2(nand_tmp_66, mux_1551_cse, fsm_output(1));
  mux_1550_nl <= MUX_s_1_2_2(mux_tmp_1549, mux_tmp_1548, fsm_output(1));
  mux_1553_cse <= MUX_s_1_2_2(mux_1552_nl, mux_1550_nl, fsm_output(4));
  or_2479_nl <= (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(0));
  mux_1546_cse <= MUX_s_1_2_2(or_2481_cse, or_2480_cse, or_2479_nl);
  mux_1564_nl <= MUX_s_1_2_2(or_tmp_611, or_tmp_330, fsm_output(3));
  attention_2_1_16_16_4_4_q_proj_re_and_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT((NOT mux_1564_nl) AND and_dcpl_581));
  or_2486_cse <= reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 OR CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd/=STD_LOGIC_VECTOR'("100"));
  or_2493_nl <= (fsm_output(5)) OR nor_tmp_285;
  mux_1580_nl <= MUX_s_1_2_2(or_2493_nl, or_2699_cse, fsm_output(3));
  or_2494_nl <= (fsm_output(6)) OR mux_1580_nl;
  mux_1581_nl <= MUX_s_1_2_2(not_tmp_253, or_2494_nl, fsm_output(7));
  attention_2_1_16_16_4_4_k_proj_re_and_1_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (mux_1581_nl OR (fsm_output(8)));
  nand_381_cse <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11")));
  or_3039_cse <= CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("00"))
      OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  APPLY_ROTARY_POS_EMB_LOOP_6_k_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c0 OR and_dcpl_726 OR APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c2
      OR APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c3 OR APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c4);
  nand_365_cse <= NOT((fsm_output(7)) AND (NOT(((RESHAPE_2D_TO_3D_LOOP_2_2_and_cse
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))) AND (fsm_output(4)))
      OR (fsm_output(5)))));
  or_2566_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10"));
  mux_1639_cse <= MUX_s_1_2_2(or_2699_cse, or_2566_nl, fsm_output(1));
  or_2576_nl <= RESHAPE_2D_TO_3D_LOOP_2_2_and_cse OR (fsm_output(2)) OR (fsm_output(3))
      OR (fsm_output(0));
  mux_1645_cse <= MUX_s_1_2_2(or_2481_cse, or_2480_cse, or_2576_nl);
  mux_1811_nl <= MUX_s_1_2_2(mux_806_cse, or_1983_cse, fsm_output(1));
  mux_1810_nl <= MUX_s_1_2_2(or_2249_cse, mux_806_cse, fsm_output(1));
  mux_1812_cse <= MUX_s_1_2_2(mux_1811_nl, mux_1810_nl, fsm_output(0));
  or_2638_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"));
  mux_1809_cse <= MUX_s_1_2_2(mux_806_cse, or_1983_cse, or_2638_nl);
  or_2671_cse <= CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01"))
      OR reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 OR (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0));
  or_2699_cse <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00"));
  and_1034_itm <= and_dcpl_732 AND and_dcpl_987;
  mux_1964_nl <= MUX_s_1_2_2(mux_1559_cse, mux_1557_cse, and_1773_cse);
  mux_1959_nl <= MUX_s_1_2_2(or_tmp_464, mux_tmp_121, or_2699_cse);
  mux_1958_nl <= MUX_s_1_2_2(mux_tmp_1549, mux_tmp_1548, fsm_output(4));
  mux_1960_nl <= MUX_s_1_2_2(mux_1959_nl, mux_1958_nl, fsm_output(1));
  mux_1954_nl <= MUX_s_1_2_2(mux_1551_cse, mux_tmp_1548, fsm_output(4));
  mux_1957_nl <= MUX_s_1_2_2(mux_1559_cse, mux_1954_nl, fsm_output(1));
  nor_540_nl <= NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("10")));
  mux_1961_nl <= MUX_s_1_2_2(mux_1960_nl, mux_1957_nl, nor_540_nl);
  mux_1962_nl <= MUX_s_1_2_2(mux_1559_cse, mux_1961_nl, and_1773_cse);
  mux_1965_nl <= MUX_s_1_2_2(mux_1964_nl, mux_1962_nl, fsm_output(0));
  or_2696_nl <= (CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11"))) OR
      (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(8));
  or_2695_nl <= (NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 OR reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      OR (fsm_output(1)) OR (NOT (fsm_output(4))))) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(8));
  mux_1948_nl <= MUX_s_1_2_2(or_2695_nl, or_2481_cse, fsm_output(2));
  mux_1949_nl <= MUX_s_1_2_2(mux_1948_nl, or_2480_cse, fsm_output(3));
  mux_1950_nl <= MUX_s_1_2_2(or_2696_nl, mux_1949_nl, fsm_output(0));
  mux_1966_itm <= MUX_s_1_2_2(mux_1965_nl, mux_1950_nl, fsm_output(7));
  and_1037_itm <= and_dcpl_743 AND and_dcpl_551 AND and_dcpl_825;
  and_1042_ssc <= and_dcpl_732 AND and_dcpl_57 AND (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(1)))
      AND and_dcpl_651;
  nor_551_nl <= NOT(CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)/=STD_LOGIC_VECTOR'("00")) OR reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 OR
      (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0))));
  mux_1982_nl <= MUX_s_1_2_2(mux_806_cse, mux_1812_cse, nor_551_nl);
  mux_1983_nl <= MUX_s_1_2_2(or_2249_cse, mux_1982_nl, and_1773_cse);
  or_2712_nl <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 OR reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"));
  mux_1976_nl <= MUX_s_1_2_2(or_1983_cse, mux_806_cse, or_2712_nl);
  mux_1975_nl <= MUX_s_1_2_2(mux_806_cse, or_1983_cse, and_1474_cse);
  mux_1977_nl <= MUX_s_1_2_2(mux_1976_nl, mux_1975_nl, fsm_output(2));
  mux_1978_nl <= MUX_s_1_2_2(mux_1977_nl, or_1983_cse, fsm_output(3));
  mux_1984_nl <= MUX_s_1_2_2(mux_1983_nl, mux_1978_nl, fsm_output(4));
  mux_1985_nl <= MUX_s_1_2_2(mux_1984_nl, or_1983_cse, fsm_output(5));
  apply_rotary_pos_emb_1_4_4_rotated_q_and_16_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (mux_1985_nl OR (fsm_output(8)));
  or_2717_cse <= (fsm_output(5)) OR mux_806_cse;
  mux_1995_nl <= MUX_s_1_2_2(mux_tmp_1993, mux_tmp_1990, fsm_output(2));
  mux_1994_nl <= MUX_s_1_2_2(mux_tmp_1993, or_2717_cse, and_1559_cse);
  nor_552_nl <= NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(0))));
  mux_1996_nl <= MUX_s_1_2_2(mux_1995_nl, mux_1994_nl, nor_552_nl);
  mux_1997_nl <= MUX_s_1_2_2(mux_tmp_1993, mux_1996_nl, fsm_output(3));
  or_2716_nl <= (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_1988_nl <= MUX_s_1_2_2(mux_806_cse, or_1983_cse, or_2716_nl);
  or_2715_nl <= (fsm_output(1)) OR (fsm_output(5));
  mux_1987_nl <= MUX_s_1_2_2(mux_806_cse, or_1983_cse, or_2715_nl);
  mux_1989_nl <= MUX_s_1_2_2(mux_1988_nl, mux_1987_nl, fsm_output(2));
  mux_1991_nl <= MUX_s_1_2_2(mux_tmp_1990, mux_1989_nl, fsm_output(0));
  mux_1992_nl <= MUX_s_1_2_2(mux_1991_nl, or_1983_cse, fsm_output(3));
  mux_1998_nl <= MUX_s_1_2_2(mux_1997_nl, mux_1992_nl, fsm_output(4));
  apply_rotary_pos_emb_1_4_4_rotated_q_and_17_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1068 OR (NOT(mux_1998_nl OR (fsm_output(8)))))) OR and_dcpl_619
      OR apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1 OR and_dcpl_1003);
  and_1762_cse <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"));
  or_2742_cse <= (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(8));
  or_2736_cse <= (fsm_output(4)) OR (fsm_output(6)) OR (NOT (fsm_output(8)));
  or_2739_cse <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("01"));
  mux_2024_cse <= MUX_s_1_2_2(or_tmp_464, mux_tmp_121, fsm_output(4));
  mux_2025_cse <= MUX_s_1_2_2(mux_2024_cse, or_2736_cse, fsm_output(5));
  mux_2032_cse <= MUX_s_1_2_2(or_2742_cse, mux_tmp_824, fsm_output(5));
  and_1055_ssc <= and_dcpl_732 AND and_dcpl_592;
  and_1059_ssc <= and_dcpl_743 AND and_dcpl_551 AND and_dcpl_835;
  or_2741_nl <= (NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd OR (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1))
      OR (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2) OR (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0))))
      OR (NOT (fsm_output(6))) OR (fsm_output(8));
  mux_2027_nl <= MUX_s_1_2_2(or_tmp_464, mux_tmp_121, or_2739_cse);
  mux_2028_nl <= MUX_s_1_2_2(or_2741_nl, mux_2027_nl, fsm_output(4));
  mux_2029_nl <= MUX_s_1_2_2(or_tmp_464, mux_2028_nl, fsm_output(0));
  mux_2030_nl <= MUX_s_1_2_2(mux_2029_nl, mux_tmp_824, fsm_output(5));
  mux_2031_nl <= MUX_s_1_2_2(mux_2030_nl, mux_2025_cse, fsm_output(1));
  mux_2033_nl <= MUX_s_1_2_2(mux_2032_cse, mux_2031_nl, and_1773_cse);
  APPLY_ROTARY_POS_EMB_LOOP_6_and_30_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (mux_2033_nl OR (fsm_output(7)));
  and_1060_itm <= and_dcpl_732 AND and_dcpl_613;
  nor_410_nl <= NOT((NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd) OR
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1)) OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2
      OR (NOT (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0))));
  mux_2036_nl <= MUX_s_1_2_2(mux_tmp_1945, mux_tmp_1943, nor_410_nl);
  apply_rotary_pos_emb_1_4_4_rotated_q_and_18_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT((NOT mux_2036_nl) AND and_dcpl_259));
  and_1062_ssc <= and_dcpl_732 AND and_dcpl_607;
  and_1626_nl <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd AND (NOT (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1)))
      AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0));
  mux_2037_nl <= MUX_s_1_2_2(mux_tmp_1945, mux_tmp_1943, and_1626_nl);
  apply_rotary_pos_emb_1_4_4_rotated_q_and_19_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT((NOT mux_2037_nl) AND and_dcpl_259));
  attention_2_1_16_16_4_4_k_proj_re_and_91_cse <= (NOT RESHAPE_2D_TO_3D_LOOP_2_2_and_cse)
      AND and_dcpl_1034;
  attention_2_1_16_16_4_4_k_proj_re_or_cse <= and_dcpl_1033 OR attention_2_1_16_16_4_4_k_proj_re_and_91_cse;
  attention_2_1_16_16_4_4_k_proj_re_or_17_cse <= (RESHAPE_2D_TO_3D_LOOP_2_2_and_cse
      AND and_dcpl_1034) OR and_dcpl_213;
  and_1771_cse <= (fsm_output(2)) AND (fsm_output(4));
  mux_2087_nl <= MUX_s_1_2_2(not_tmp_874, or_tmp_1132, fsm_output(7));
  mux_2086_nl <= MUX_s_1_2_2(not_tmp_874, or_tmp_1218, fsm_output(7));
  mux_2088_nl <= MUX_s_1_2_2(mux_2087_nl, mux_2086_nl, reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  nor_1228_ssc <= NOT(mux_2088_nl OR (fsm_output(8)));
  nand_357_nl <= NOT((fsm_output(6)) AND mux_tmp_1489);
  mux_1542_nl <= MUX_s_1_2_2(nand_357_nl, or_tmp_1132, fsm_output(7));
  attention_2_1_16_16_4_4_q_proj_and_5_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (mux_1542_nl OR (fsm_output(8)) OR and_dcpl_626);
  or_2792_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"));
  or_2797_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"));
  mux_2092_cse <= MUX_s_1_2_2(or_2457_cse, or_1197_cse, fsm_output(4));
  or_2799_nl <= (NOT (fsm_output(0))) OR (fsm_output(1)) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (fsm_output(8));
  mux_2097_nl <= MUX_s_1_2_2(or_2460_cse, or_tmp_1643, or_1732_cse);
  mux_2098_nl <= MUX_s_1_2_2(or_2799_nl, mux_2097_nl, fsm_output(3));
  mux_2096_nl <= MUX_s_1_2_2(mux_1522_cse, or_1197_cse, or_2797_cse);
  mux_2099_nl <= MUX_s_1_2_2(mux_2098_nl, mux_2096_nl, fsm_output(5));
  mux_2093_nl <= MUX_s_1_2_2(mux_2092_cse, or_tmp_1643, or_2792_cse);
  mux_2094_nl <= MUX_s_1_2_2(or_2460_cse, mux_2093_nl, fsm_output(3));
  or_2787_nl <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(4));
  mux_2090_nl <= MUX_s_1_2_2(mux_1522_cse, or_1197_cse, or_2787_nl);
  or_2786_nl <= ((fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(4))) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100"));
  mux_2091_nl <= MUX_s_1_2_2(mux_2090_nl, or_2786_nl, fsm_output(3));
  mux_2095_nl <= MUX_s_1_2_2(mux_2094_nl, mux_2091_nl, fsm_output(5));
  mux_2100_ssc <= MUX_s_1_2_2(mux_2099_nl, mux_2095_nl, fsm_output(2));
  APPLY_ROTARY_POS_EMB_LOOP_6_and_28_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (and_dcpl_888 OR and_dcpl_257 OR and_dcpl_1073 OR and_dcpl_240 OR and_dcpl_207
      OR and_dcpl_847 OR and_dcpl_583);
  APPLY_ROTARY_POS_EMB_LOOP_6_and_31_cse <= APPLY_ROTARY_POS_EMB_LOOP_6_and_28_cse
      AND (NOT and_dcpl_725);
  nand_283_nl <= NOT((fsm_output(6)) AND mux_tmp_1421);
  mux_2102_nl <= MUX_s_1_2_2(nand_283_nl, or_tmp_1218, fsm_output(7));
  attention_2_1_16_16_4_4_q_proj_re_and_29_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (mux_2102_nl OR (fsm_output(8)));
  mux_2103_nl <= MUX_s_1_2_2((NOT or_tmp_728), or_tmp_762, fsm_output(5));
  mux_2104_nl <= MUX_s_1_2_2(mux_tmp_91, mux_2103_nl, fsm_output(3));
  attention_2_1_16_16_4_4_k_proj_re_and_65_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT((NOT mux_2104_nl) AND and_dcpl_259));
  attention_2_1_16_16_4_4_v_proj_re_and_32_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT(((and_1638_cse OR (fsm_output(4))) XOR (fsm_output(5))) AND and_dcpl_259));
  LINEAR_FORWARD_NO_MUL_LOOP_2_and_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT((NOT (fsm_output(2))) OR (fsm_output(4)) OR (fsm_output(8)) OR nand_197_cse
      OR or_dcpl_1134 OR or_1983_cse));
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_and_29_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (and_dcpl_257 OR and_dcpl_410 OR and_dcpl_240 OR and_dcpl_1034 OR and_dcpl_207
      OR and_dcpl_213 OR and_dcpl_583 OR and_dcpl_265);
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse <= and_dcpl_410 OR attention_2_1_16_16_4_4_k_proj_re_and_91_cse;
  nand_285_nl <= NOT((fsm_output(6)) AND mux_tmp_857);
  or_2828_nl <= (fsm_output(5)) OR nor_tmp_282;
  mux_2107_nl <= MUX_s_1_2_2(or_2828_nl, or_2699_cse, fsm_output(3));
  or_3153_nl <= (fsm_output(6)) OR mux_2107_nl;
  mux_2108_nl <= MUX_s_1_2_2(nand_285_nl, or_3153_nl, fsm_output(7));
  attention_2_1_16_16_4_4_v_proj_re_and_95_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (mux_2108_nl OR (fsm_output(8)));
  mux_2109_nl <= MUX_s_1_2_2(nor_717_cse, or_3137_cse, fsm_output(3));
  attention_2_1_16_16_4_4_v_proj_and_30_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT((NOT(mux_2109_nl OR (fsm_output(8)))) AND and_dcpl_1145));
  GEMM_3D_FLOAT_LOOP_3_1_mux_4_nl <= MUX_s_1_2_2((NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1),
      (NOT or_dcpl_1155), and_dcpl_1154);
  mux_2124_nl <= MUX_s_1_2_2(nand_tmp_99, or_tmp_1664, or_270_cse);
  mux_2123_nl <= MUX_s_1_2_2(mux_tmp_2116, or_tmp_1671, fsm_output(2));
  mux_2125_nl <= MUX_s_1_2_2(mux_2124_nl, mux_2123_nl, fsm_output(3));
  mux_2126_nl <= MUX_s_1_2_2(mux_2125_nl, mux_tmp_2121, fsm_output(1));
  or_2840_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 5)/=STD_LOGIC_VECTOR'("1000"));
  mux_2114_nl <= MUX_s_1_2_2(or_tmp_1664, or_2840_nl, and_1771_cse);
  mux_2120_nl <= MUX_s_1_2_2(mux_tmp_2119, mux_2114_nl, fsm_output(3));
  mux_2122_nl <= MUX_s_1_2_2(mux_tmp_2121, mux_2120_nl, fsm_output(1));
  mux_2127_nl <= MUX_s_1_2_2(mux_2126_nl, mux_2122_nl, fsm_output(0));
  GEMM_3D_FLOAT_LOOP_3_1_and_44_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((GEMM_3D_FLOAT_LOOP_3_1_mux_4_nl AND mux_2127_nl) OR and_dcpl_1152 OR
      and_dcpl_222);
  mux_2128_nl <= MUX_s_1_2_2(or_3167_cse, or_1907_cse, fsm_output(0));
  attention_2_1_16_16_4_4_q_embed_and_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT((NOT mux_2128_nl) AND and_dcpl_201 AND and_dcpl_199));
  and_1782_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111"));
  nor_1239_cse <= NOT((fsm_output(5)) OR and_1782_cse OR (fsm_output(6)) OR (NOT
      (fsm_output(8))));
  nor_593_cse <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")));
  nor_1240_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_1241_nl <= NOT((NOT((fsm_output(4)) OR (fsm_output(6)))) OR (fsm_output(8)));
  mux_2155_nl <= MUX_s_1_2_2(nor_1240_nl, nor_1241_nl, and_1474_cse);
  nor_1242_nl <= NOT((NOT((NOT((fsm_output(1)) OR (fsm_output(0)) OR (NOT (fsm_output(4)))))
      OR (fsm_output(6)))) OR (fsm_output(8)));
  mux_2156_nl <= MUX_s_1_2_2(mux_2155_nl, nor_1242_nl, fsm_output(2));
  nor_1243_nl <= NOT((NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_1244_nl <= NOT((NOT((NOT((fsm_output(0)) OR (z_out_5(2)))) OR (fsm_output(4))))
      OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_2154_nl <= MUX_s_1_2_2(nor_1243_nl, nor_1244_nl, nor_593_cse);
  mux_2157_cse <= MUX_s_1_2_2(mux_2156_nl, mux_2154_nl, fsm_output(3));
  attention_2_1_16_16_4_4_attn_weights_and_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT(and_dcpl_185 AND or_1732_cse AND and_dcpl_190));
  GEMM_3D_FLOAT_LOOP_3_and_36_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT((or_1732_cse XOR (fsm_output(2))) AND and_dcpl_61 AND and_dcpl_190));
  attention_2_1_16_16_4_4_attn_weights_and_52_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT(and_dcpl_61 AND (NOT (fsm_output(2))) AND (fsm_output(5)) AND and_dcpl_1141));
  attention_2_1_16_16_4_4_attn_weights_and_48_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT and_dcpl_1195);
  mux_1543_nl <= MUX_s_1_2_2((NOT (fsm_output(2))), (fsm_output(2)), fsm_output(1));
  mux_2237_nl <= MUX_s_1_2_2(or_3167_cse, mux_1543_nl, fsm_output(0));
  attention_2_1_16_16_4_4_attn_weights_and_12_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT((NOT mux_2237_nl) AND and_dcpl_61 AND and_dcpl_293));
  attention_2_1_16_16_4_4_attn_weights_and_24_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT and_dcpl_304);
  GEMM_3D_FLOAT_LOOP_3_1_and_46_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT((NOT(mux_tmp_1440 OR (fsm_output(8)))) AND nor_646_cse AND and_dcpl_148));
  mux_2249_nl <= MUX_s_1_2_2((NOT nor_tmp_285), or_tmp_861, fsm_output(5));
  mux_2250_nl <= MUX_s_1_2_2(mux_2249_nl, or_tmp_682, fsm_output(3));
  attention_abs_4_qelse_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT((NOT mux_2250_nl) AND and_dcpl_258 AND (fsm_output(7))));
  compute_sqrt_1_guess_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((and_dcpl_362 AND and_dcpl_221) OR and_dcpl_292);
  attention_2_1_16_16_4_4_quantized_final_output_and_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1158 OR (NOT mux_2256_itm))) OR mux_tmp_2252);
  RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse <= (NOT QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1)
      AND and_dcpl_1154;
  RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse <= QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1
      AND and_dcpl_1154;
  attention_2_1_16_16_4_4_quantized_final_output_and_8_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1166 OR (NOT mux_2256_itm))) OR mux_tmp_2252);
  attention_2_1_16_16_4_4_quantized_final_output_and_16_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1164 OR (NOT mux_2256_itm))) OR mux_tmp_2252);
  attention_2_1_16_16_4_4_quantized_final_output_and_24_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1161 OR (NOT mux_2256_itm))) OR mux_tmp_2252);
  attention_2_1_16_16_4_4_quantized_final_output_and_32_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1159 OR (NOT mux_2256_itm))) OR mux_tmp_2252);
  attention_2_1_16_16_4_4_quantized_final_output_and_40_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1156 OR (NOT mux_2256_itm))) OR mux_tmp_2252);
  attention_2_1_16_16_4_4_quantized_final_output_and_48_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1160 OR (NOT mux_2256_itm))) OR mux_tmp_2252);
  attention_2_1_16_16_4_4_quantized_final_output_and_56_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1162 OR (NOT mux_2256_itm))) OR mux_tmp_2252);
  attention_2_1_16_16_4_4_quantized_final_output_and_64_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1165 OR (NOT mux_2256_itm))) OR mux_tmp_2252);
  attention_2_1_16_16_4_4_quantized_final_output_and_72_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1167 OR (NOT mux_2256_itm))) OR mux_tmp_2252);
  attention_2_1_16_16_4_4_quantized_final_output_and_80_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1169 OR (NOT mux_2256_itm))) OR mux_tmp_2252);
  attention_2_1_16_16_4_4_quantized_final_output_and_88_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1141 OR (NOT mux_2256_itm))) OR mux_tmp_2252);
  attention_2_1_16_16_4_4_quantized_final_output_and_96_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1170 OR (NOT mux_2256_itm))) OR mux_tmp_2252);
  attention_2_1_16_16_4_4_quantized_final_output_and_104_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND ((NOT(or_dcpl_1168 OR (NOT mux_2256_itm))) OR mux_tmp_2252);
  mux_2257_nl <= MUX_s_1_2_2(or_dcpl_1050, nor_tmp_329, fsm_output(5));
  mux_2258_nl <= MUX_s_1_2_2((fsm_output(5)), (NOT mux_2257_nl), fsm_output(3));
  attention_2_1_16_16_4_4_quantized_final_output_and_112_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (NOT(mux_2258_nl AND and_dcpl_413));
  attention_2_1_16_16_4_4_v_proj_re_and_63_cse <= (NOT or_dcpl_1141) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_65_cse <= (NOT or_dcpl_1170) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_67_cse <= (NOT or_dcpl_1169) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_69_cse <= (NOT or_dcpl_1168) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_71_cse <= (NOT or_dcpl_1167) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_73_cse <= (NOT or_dcpl_1166) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_75_cse <= (NOT or_dcpl_1165) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_77_cse <= (NOT or_dcpl_1164) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_79_cse <= (NOT or_dcpl_1162) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_81_cse <= (NOT or_dcpl_1161) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_83_cse <= (NOT or_dcpl_1160) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_85_cse <= (NOT or_dcpl_1159) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_87_cse <= (NOT or_dcpl_1158) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_89_cse <= (NOT or_dcpl_1156) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_91_cse <= (NOT or_dcpl_1155) AND and_dcpl_1225;
  attention_2_1_16_16_4_4_v_proj_re_and_93_cse <= (NOT or_dcpl_1152) AND and_dcpl_1225;
  output_and_16_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT(((and_1771_cse
      AND (fsm_output(1)) AND (fsm_output(3))) XOR (fsm_output(5))) AND and_dcpl_413));
  output_and_64_cse <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT
      and_dcpl_1232);
  or_1659_nl <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd OR (NOT GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva);
  attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2_mx1 <= MUX_v_40_2_2(acc_3_cse_40_1,
      attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3, or_1659_nl);
  nand_298_nl <= NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd AND LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0);
  attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2_mx1 <= MUX_v_40_2_2(acc_3_cse_40_1,
      attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3, nand_298_nl);
  or_1661_nl <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd OR (NOT GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva);
  attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2_mx1 <= MUX_v_40_2_2(acc_3_cse_40_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2, or_1661_nl);
  nand_299_nl <= NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd AND reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2_mx1 <= MUX_v_40_2_2(acc_3_cse_40_1,
      attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3, nand_299_nl);
  or_1663_nl <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd OR (NOT GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva);
  attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2_mx1 <= MUX_v_40_2_2(acc_3_cse_40_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2, or_1663_nl);
  nand_300_nl <= NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd AND GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva);
  attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2_mx1 <= MUX_v_40_2_2(acc_3_cse_40_1,
      attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3, nand_300_nl);
  or_1665_nl <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd OR (NOT GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva);
  attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2_mx1 <= MUX_v_40_2_2(acc_3_cse_40_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2, or_1665_nl);
  nand_301_nl <= NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd AND GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva);
  attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2_mx1 <= MUX_v_40_2_2(acc_3_cse_40_1,
      attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3, nand_301_nl);
  or_1667_ssc <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd OR (NOT GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva);
  attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_39 <= MUX_s_1_2_2((acc_3_cse_40_1(39)),
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd, or_1667_ssc);
  attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_38_0 <= MUX_v_39_2_2((acc_3_cse_40_1(38
      DOWNTO 0)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1, or_1667_ssc);
  or_1669_nl <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd OR (NOT GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva);
  attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2_mx1 <= MUX_v_40_2_2(acc_3_cse_40_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2, or_1669_nl);
  or_1671_nl <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd OR (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2_mx1 <= MUX_v_40_2_2(acc_3_cse_40_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2, or_1671_nl);
  attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2_mx1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva);
  attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2_mx1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_1,
      acc_3_cse_40_1, reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2_mx1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva);
  attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2_mx1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_1,
      acc_3_cse_40_1, LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0);
  attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2_mx1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva);
  attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2_mx1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva);
  attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2_mx1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva);
  attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2_mx1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva);
  attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2_mx1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva);
  attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2_mx1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva);
  attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2_mx1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva);
  attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2_mx1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_sva);
  attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1, or_dcpl_980);
  attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1, or_dcpl_983);
  attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1, or_dcpl_985);
  attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1, or_dcpl_989);
  attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1, or_dcpl_990);
  attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1, or_dcpl_993);
  attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1, or_dcpl_998);
  attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3, or_dcpl_980);
  attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3, or_dcpl_983);
  attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3, or_dcpl_985);
  attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3, or_dcpl_987);
  attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2, or_dcpl_988);
  attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3, or_dcpl_989);
  and_1455_cse <= (((fsm_output(4)) AND (fsm_output(6))) OR (fsm_output(7))) AND
      (fsm_output(8));
  nor_176_cse <= NOT((fsm_output(1)) OR (NOT (fsm_output(4))));
  attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2, or_dcpl_990);
  attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2, or_dcpl_993);
  attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2, or_dcpl_996);
  attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2, or_dcpl_998);
  attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1, or_dcpl_1000);
  attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_39_16, or_dcpl_1002);
  attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_15_0, or_dcpl_1002);
  attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_39_16, or_dcpl_1004);
  attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_15_0, or_dcpl_1004);
  attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_39_16, or_dcpl_1006);
  attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_15_0, or_dcpl_1006);
  attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16, or_dcpl_1008);
  attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_15_0, or_dcpl_1008);
  attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_39_16, or_dcpl_1009);
  attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_15_0, or_dcpl_1009);
  attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16, or_dcpl_1010);
  attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_39_16, or_dcpl_1011);
  attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_15_0, or_dcpl_1011);
  attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16, or_dcpl_1012);
  attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_39_16, or_dcpl_1013);
  attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0, or_dcpl_1013);
  attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16, or_dcpl_1014);
  attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_39_16, or_dcpl_1015);
  attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_15_0, or_dcpl_1015);
  attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16, or_dcpl_1016);
  attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_39_16, or_dcpl_1017);
  attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_15_0, or_dcpl_1017);
  attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16, or_dcpl_1018);
  attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16, or_dcpl_1019);
  attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_15_0, or_dcpl_1019);
  apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2, or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2, or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w0 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2, or_dcpl_1023);
  mux_502_cse <= MUX_s_1_2_2(or_2456_cse, (fsm_output(8)), fsm_output(7));
  apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w3 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2, or_dcpl_1025);
  apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2_mx0w1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16_mx0w1 <= MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1,
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 <= MUX_v_8_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm,
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16_mx0w1 <= MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_39_16, or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_13 <= MUX_v_3_2_2((APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm(7
      DOWNTO 5)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd,
      or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_12_8 <= MUX_v_5_2_2((APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm(4
      DOWNTO 0)), (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1(12
      DOWNTO 8)), or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1(7)), or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1(6)), or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1(5)), or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1(4)), or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1(3)), or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1(2)), or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1(1)), or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1(0)), or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16_mx0w1 <= MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_39_16, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 <= MUX_v_8_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_15_8, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_7, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_6, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_5, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_4, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_3, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_2, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_1, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_0, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 <= MUX_v_8_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0, or_dcpl_1023);
  apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16_mx0w1 <= MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16, or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 <= MUX_v_8_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd, or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7, or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6, or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5, or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4, or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3, or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2, or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1, or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0, or_dcpl_1021);
  apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16_mx0w1 <= MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_39_16, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 <= MUX_v_8_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1, or_dcpl_1024);
  apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0 <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0, or_dcpl_1024);
  attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out(15
      DOWNTO 8)), attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_15_8, or_dcpl_1028);
  attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out(7)),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7, or_dcpl_1028);
  attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out(6)),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6, or_dcpl_1028);
  attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out(5)),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5, or_dcpl_1028);
  attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out(4)),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4, or_dcpl_1028);
  attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out(3)),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3, or_dcpl_1028);
  attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out(2)),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2, or_dcpl_1028);
  attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out(1)),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1, or_dcpl_1028);
  attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out(0)),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0, or_dcpl_1028);
  attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out(15
      DOWNTO 8)), attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_15_8, or_dcpl_1030);
  attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out(7)),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7, or_dcpl_1030);
  attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out(6)),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6, or_dcpl_1030);
  attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out(5)),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5, or_dcpl_1030);
  attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out(4)),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4, or_dcpl_1030);
  attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out(3)),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3, or_dcpl_1030);
  attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out(2)),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2, or_dcpl_1030);
  attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out(1)),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1, or_dcpl_1030);
  attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out(0)),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0, or_dcpl_1030);
  attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out(15
      DOWNTO 8)), attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_15_8, or_dcpl_1031);
  attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out(7)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7, or_dcpl_1031);
  attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out(6)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6, or_dcpl_1031);
  attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out(5)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5, or_dcpl_1031);
  attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out(4)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4, or_dcpl_1031);
  attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out(3)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3, or_dcpl_1031);
  attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out(2)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2, or_dcpl_1031);
  attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out(1)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1, or_dcpl_1031);
  attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out(0)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0, or_dcpl_1031);
  attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out(15
      DOWNTO 8)), attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_15_8, or_dcpl_1033);
  attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out(7)),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7, or_dcpl_1033);
  attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out(6)),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6, or_dcpl_1033);
  attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out(5)),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5, or_dcpl_1033);
  attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out(4)),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4, or_dcpl_1033);
  attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out(3)),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3, or_dcpl_1033);
  attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out(2)),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2, or_dcpl_1033);
  attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out(1)),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1, or_dcpl_1033);
  attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out(0)),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0, or_dcpl_1033);
  attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out(15
      DOWNTO 8)), attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_15_8, or_dcpl_1035);
  attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out(7)),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7, or_dcpl_1035);
  attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out(6)),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6, or_dcpl_1035);
  attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out(5)),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5, or_dcpl_1035);
  attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out(4)),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4, or_dcpl_1035);
  attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out(3)),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3, or_dcpl_1035);
  attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out(2)),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2, or_dcpl_1035);
  attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out(1)),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1, or_dcpl_1035);
  attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out(0)),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0, or_dcpl_1035);
  attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out(15
      DOWNTO 8)), attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_15_8, or_dcpl_1037);
  attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out(7)),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7, or_dcpl_1037);
  attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out(6)),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6, or_dcpl_1037);
  attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out(5)),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5, or_dcpl_1037);
  attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out(4)),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4, or_dcpl_1037);
  attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out(3)),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3, or_dcpl_1037);
  attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out(2)),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2, or_dcpl_1037);
  attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out(1)),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1, or_dcpl_1037);
  attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out(0)),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0, or_dcpl_1037);
  attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out(15
      DOWNTO 8)), attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_8, or_dcpl_1038);
  attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out(7)),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd, or_dcpl_1038);
  attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out(6)),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_1, or_dcpl_1038);
  attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out(5)),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_2, or_dcpl_1038);
  attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out(4)),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_3, or_dcpl_1038);
  attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out(3)),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_4, or_dcpl_1038);
  attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out(2)),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_5, or_dcpl_1038);
  attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out(1)),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_6, or_dcpl_1038);
  attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out(0)),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_7, or_dcpl_1038);
  attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out(15
      DOWNTO 8)), attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_15_8, or_dcpl_1039);
  attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out(7)),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_7, or_dcpl_1039);
  attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out(6)),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_6, or_dcpl_1039);
  attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out(5)),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_5, or_dcpl_1039);
  attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out(4)),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_4, or_dcpl_1039);
  attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out(3)),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_3, or_dcpl_1039);
  attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out(2)),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_2, or_dcpl_1039);
  attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out(1)),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_1, or_dcpl_1039);
  attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out(0)),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_0, or_dcpl_1039);
  attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out(15
      DOWNTO 8)), attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_15_8, or_dcpl_1041);
  attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out(7)),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7, or_dcpl_1041);
  attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out(6)),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6, or_dcpl_1041);
  attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out(5)),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5, or_dcpl_1041);
  attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out(4)),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4, or_dcpl_1041);
  attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out(3)),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3, or_dcpl_1041);
  attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out(2)),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2, or_dcpl_1041);
  attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out(1)),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1, or_dcpl_1041);
  attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out(0)),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0, or_dcpl_1041);
  attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(z_out, attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_15_0,
      or_dcpl_1042);
  attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out(15
      DOWNTO 8)), attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_15_8, or_dcpl_1043);
  attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out(7)),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7, or_dcpl_1043);
  attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out(6)),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6, or_dcpl_1043);
  attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out(5)),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5, or_dcpl_1043);
  attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out(4)),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4, or_dcpl_1043);
  attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out(3)),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3, or_dcpl_1043);
  attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out(2)),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2, or_dcpl_1043);
  attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out(1)),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1, or_dcpl_1043);
  attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out(0)),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0, or_dcpl_1043);
  attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(z_out, attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_15_0,
      or_dcpl_1044);
  attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out(15
      DOWNTO 8)), attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_15_8, or_dcpl_1045);
  attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out(7)),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7, or_dcpl_1045);
  attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out(6)),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6, or_dcpl_1045);
  attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out(5)),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5, or_dcpl_1045);
  attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out(4)),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4, or_dcpl_1045);
  attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out(3)),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3, or_dcpl_1045);
  attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out(2)),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2, or_dcpl_1045);
  attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out(1)),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1, or_dcpl_1045);
  attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out(0)),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0, or_dcpl_1045);
  attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out(15
      DOWNTO 8)), attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_15_8, or_dcpl_1046);
  attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out(7)),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7, or_dcpl_1046);
  attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out(6)),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6, or_dcpl_1046);
  attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out(5)),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5, or_dcpl_1046);
  attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out(4)),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4, or_dcpl_1046);
  attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out(3)),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3, or_dcpl_1046);
  attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out(2)),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2, or_dcpl_1046);
  attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out(1)),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1, or_dcpl_1046);
  attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out(0)),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0, or_dcpl_1046);
  attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16, or_dcpl_1002);
  attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out_1(15
      DOWNTO 8)), apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_15_8, or_dcpl_1002);
  attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out_1(7)),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_7, or_dcpl_1002);
  attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out_1(6)),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_6, or_dcpl_1002);
  attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out_1(5)),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_5, or_dcpl_1002);
  attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out_1(4)),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_4, or_dcpl_1002);
  attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out_1(3)),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_3, or_dcpl_1002);
  attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out_1(2)),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_2, or_dcpl_1002);
  attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out_1(1)),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_1, or_dcpl_1002);
  attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out_1(0)),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_0, or_dcpl_1002);
  attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_39_16, or_dcpl_1004);
  attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0, or_dcpl_1004);
  attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_39_16, or_dcpl_1006);
  attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_15_13 <= MUX_v_3_2_2((z_out_1(15
      DOWNTO 13)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd,
      or_dcpl_1006);
  attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0 <= MUX_v_13_2_2((z_out_1(12
      DOWNTO 0)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1,
      or_dcpl_1006);
  attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_39_16, or_dcpl_1008);
  attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_15_0, or_dcpl_1008);
  attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_39_16, or_dcpl_1009);
  attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(z_out_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0, or_dcpl_1009);
  attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_39_16, or_dcpl_1010);
  attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_15_0, or_dcpl_1010);
  attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48, or_dcpl_1011);
  attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_39_16, or_dcpl_1012);
  attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0, or_dcpl_1012);
  attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_39_16, or_dcpl_1013);
  attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out_1(15
      DOWNTO 8)), APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8, or_dcpl_1013);
  attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out_1(7)),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7, or_dcpl_1013);
  attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out_1(6)),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6, or_dcpl_1013);
  attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out_1(5)),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5, or_dcpl_1013);
  attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out_1(4)),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4, or_dcpl_1013);
  attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out_1(3)),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3, or_dcpl_1013);
  attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out_1(2)),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2, or_dcpl_1013);
  attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out_1(1)),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1, or_dcpl_1013);
  attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out_1(0)),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0, or_dcpl_1013);
  attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_39_16, or_dcpl_1014);
  attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_15_0, or_dcpl_1014);
  attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16, or_dcpl_1015);
  attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out_1(15
      DOWNTO 8)), reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd, or_dcpl_1015);
  attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out_1(7)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7, or_dcpl_1015);
  attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out_1(6)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6, or_dcpl_1015);
  attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out_1(5)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5, or_dcpl_1015);
  attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out_1(4)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4, or_dcpl_1015);
  attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out_1(3)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3, or_dcpl_1015);
  attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out_1(2)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2, or_dcpl_1015);
  attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out_1(1)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1, or_dcpl_1015);
  attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out_1(0)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0, or_dcpl_1015);
  attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_39_16, or_dcpl_1016);
  attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_15_0, or_dcpl_1016);
  attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_15_8 <= MUX_v_8_2_2((z_out_1(15
      DOWNTO 8)), reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd, or_dcpl_1017);
  attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_7 <= MUX_s_1_2_2((z_out_1(7)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7, or_dcpl_1017);
  attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_6 <= MUX_s_1_2_2((z_out_1(6)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6, or_dcpl_1017);
  attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_5 <= MUX_s_1_2_2((z_out_1(5)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5, or_dcpl_1017);
  attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_4 <= MUX_s_1_2_2((z_out_1(4)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4, or_dcpl_1017);
  attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_3 <= MUX_s_1_2_2((z_out_1(3)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3, or_dcpl_1017);
  attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_2 <= MUX_s_1_2_2((z_out_1(2)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2, or_dcpl_1017);
  attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_1 <= MUX_s_1_2_2((z_out_1(1)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1, or_dcpl_1017);
  attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_0 <= MUX_s_1_2_2((z_out_1(0)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0, or_dcpl_1017);
  attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_39_16, or_dcpl_1018);
  attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_15_0, or_dcpl_1018);
  attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16_mx0w1 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_39_16, or_dcpl_1019);
  attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0_mx0w1 <= MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_15_0, or_dcpl_1019);
  nor_749_cse <= NOT((fsm_output(2)) OR (fsm_output(0)));
  or_76_cse <= reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 OR reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd;
  or_130_cse <= (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1) OR reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd;
  drf_output_sdt_2_sva_15_0_mx0w0 <= MUX_v_16_16_2(attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0,
      (APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8 & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6 & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4 & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2 & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0), attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_15_0,
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0, attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_15_0,
      attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_15_0, attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_15_0,
      attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0, attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_15_0,
      attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_15_0, (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd
      & reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_15_8
      & apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_7 & apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_6
      & apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_5 & apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_4
      & apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_3 & apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_2
      & apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_1 & apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_0),
      attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0, attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_15_0,
      attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_15_0, attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  drf_output_sdt_3_sva_15_0_mx0w3 <= MUX_v_16_16_2(attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0,
      (APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8 & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6 & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4 & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2 & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0), apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0,
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0, attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0, reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2);
  SOFTMAX_LOOP_5_mux_12_psp_mx0w0 <= MUX_v_40_12_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_5,
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_5, attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_5,
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_5, attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_4,
      attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_4, attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_4,
      attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_4, attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_4,
      attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_4, attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_4,
      attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_4, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_conc_1_mut_71_48_mx0w0 <= MUX_v_24_16_2(attention_2_1_16_16_4_4_v_proj_re_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_3_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_4_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_5_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_6_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_7_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_8_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_9_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_10_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_12_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_13_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_14_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_15_sva_1_39_16, reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  LINEAR_FORWARD_NO_MUL_LOOP_2_3_conc_1_mut_71_48_mx0w3 <= MUX_v_24_16_2(output_0_0_sva_1_39_16,
      output_0_1_sva_1_39_16, output_0_2_sva_1_39_16, output_0_3_sva_1_39_16, output_0_4_sva_1_39_16,
      output_0_5_sva_1_39_16, output_0_6_sva_1_39_16, output_0_7_sva_1_39_16, output_0_8_sva_1_39_16,
      output_0_9_sva_1_39_16, output_0_10_sva_1_39_16, output_0_11_sva_1_39_16, output_0_12_sva_1_39_16,
      output_0_13_sva_1_39_16, output_0_14_sva_1_39_16, output_0_15_sva_1_39_16,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2);
  compute_sqrt_1_for_acc_1_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_SIGNED(SIGNED(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4
      & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0 & compute_sqrt_1_guess_sva_34
      & compute_sqrt_1_guess_sva_33_0), 40), 41) + CONV_SIGNED(CONV_SIGNED(SIGNED(APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm(39
      DOWNTO 0)), 40), 41), 41));
  compute_sqrt_1_for_acc_1_itm_40_1_1 <= compute_sqrt_1_for_acc_1_nl(40 DOWNTO 1);
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'(
      SIGNED(GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm) * SIGNED'( "0100101101010110010011")),
      61));
  or_1860_nl <= reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 OR (CM_LOOP_3_acc_tmp(0));
  attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx1 <= MUX_v_40_2_2(CM_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_ctmp_sva_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_3, or_1860_nl);
  attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx2 <= MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z(39
      DOWNTO 0)), attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_5, or_dcpl_1063);
  attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_39 <= reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      AND attention_max_attn_fixed_t_1_acc_1_itm_40_1;
  attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_38_0 <= MUX_v_39_2_2(STD_LOGIC_VECTOR'("000000000000000000000000000000000000000"),
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1, attention_max_attn_fixed_t_1_acc_1_itm_40_1);
  compute_sqrt_for_acc_1_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_SIGNED(SIGNED(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4
      & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0 & compute_sqrt_guess_sva_34
      & compute_sqrt_guess_sva_33_0), 40), 41) + CONV_SIGNED(CONV_SIGNED(SIGNED(APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm(39
      DOWNTO 0)), 40), 41), 41));
  compute_sqrt_for_acc_1_itm_40_1_1 <= compute_sqrt_for_acc_1_nl(40 DOWNTO 1);
  attention_abs_1_qr_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(NOT
      (input_0_0_sva_2(38 DOWNTO 0))), 39), 40) + SIGNED'( "0000000000000000000000000000000000000001"),
      40));
  softmax_1_4_3_sum_sva_2 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1) + SIGNED(SOFTMAX_LOOP_4_acc_3_cse_sva_1),
      40));
  attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx2 <= MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z(39
      DOWNTO 0)), attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_5, or_dcpl_1076);
  attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx1 <= MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z(39
      DOWNTO 0)), attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_4, or_dcpl_1081);
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2),
      4), 5) + SIGNED'( "00001"), 5));
  RMS_NORM_LOOP_2_2_acc_1_tmp <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
      & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1), 4), 5) + SIGNED'( "00001"), 5));
  attention_abs_qr_35_0_lpi_1_dfm_mx0w0 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(NOT
      (operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1(34
      DOWNTO 0))), 35), 36) + SIGNED'( "000000000000000000000000000000000001"), 36));
  attention_abs_qr_35_0_lpi_1_dfm_mx1_35 <= (attention_abs_qr_35_0_lpi_1_dfm_mx0w0(35))
      AND (operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1(35));
  attention_abs_qr_35_0_lpi_1_dfm_mx1_34_1 <= MUX_v_34_2_2((operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1(34
      DOWNTO 1)), (attention_abs_qr_35_0_lpi_1_dfm_mx0w0(34 DOWNTO 1)), operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1(35));
  operator_40_24_true_AC_TRN_AC_WRAP_and_1_nl <= reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd
      AND reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1
      <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd
      & (reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(38 DOWNTO 4))) + CONV_SIGNED(CONV_UNSIGNED(operator_40_24_true_AC_TRN_AC_WRAP_and_1_nl,
      1), 36), 36));
  QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_dfm_1_38_0_1 <= MUX1HOT_v_39_5_2((input_0_0_sva_2(38
      DOWNTO 0)), reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1, QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_38_0,
      (RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva(38 DOWNTO 0)), attention_abs_3_qr_sva_38_0,
      STD_LOGIC_VECTOR'( RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_nor_1_ssc_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & RMS_NORM_LOOP_2_and_29_ssc & RMS_NORM_LOOP_2_and_33_ssc_1 & RMS_NORM_LOOP_2_and_34_ssc));
  RMS_NORM_LOOP_2_2_unequal_tmp_mx0w0 <= NOT(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4
      AND CONV_SL_1_1(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0=STD_LOGIC_VECTOR'("1111")));
  TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(z_out_11(2
      DOWNTO 1)), 2), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1), 2), 3), 3));
  GEMM_3D_FLOAT_LOOP_3_acc_6_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(z_out_11(2
      DOWNTO 1)), 2), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1), 2), 3), 3));
  attention_abs_2_mux_2 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(NOT
      (RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva(38 DOWNTO 0))), 39),
      40) + SIGNED'( "0000000000000000000000000000000000000001"), 40));
  QUANTIZE_ACTIVATION_LOOP_2_attention_abs_2_nand_nl <= NOT((attention_abs_2_mux_2(39))
      AND (RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva(39)));
  attention_abs_2_mux_3_nl <= MUX_v_39_2_2((RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva(38
      DOWNTO 0)), (attention_abs_2_mux_2(38 DOWNTO 0)), RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva(39));
  QUANTIZE_ACTIVATION_LOOP_2_acc_4_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_SIGNED(SIGNED(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      & QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_38_0), 40), 41) + CONV_UNSIGNED(CONV_SIGNED(SIGNED(QUANTIZE_ACTIVATION_LOOP_2_attention_abs_2_nand_nl
      & (NOT attention_abs_2_mux_3_nl)), 40), 41) + UNSIGNED'( "00000000000000000000000000000000000000001"),
      41));
  QUANTIZE_ACTIVATION_LOOP_2_acc_4_itm_40_1 <= QUANTIZE_ACTIVATION_LOOP_2_acc_4_nl(40);
  RMS_NORM_LOOP_2_and_29_ssc_1 <= (NOT QUANTIZE_ACTIVATION_LOOP_2_acc_4_itm_40_1)
      AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  RMS_NORM_LOOP_2_and_34_ssc_1 <= (RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva(39))
      AND RMS_NORM_LOOP_2_and_30_m1c_1;
  RMS_NORM_LOOP_2_and_30_m1c_1 <= QUANTIZE_ACTIVATION_LOOP_2_acc_4_itm_40_1 AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  RMS_NORM_LOOP_2_2_and_32_ssc_mx0w3 <= (attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_2_mx0(39))
      AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_nor_1_ssc_1 <= NOT((input_0_0_sva_2(39)) OR reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  RMS_NORM_LOOP_2_and_33_ssc_1 <= (NOT (RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva(39)))
      AND RMS_NORM_LOOP_2_and_30_m1c;
  QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_dfm_1_38_0_mx0w1 <= MUX1HOT_v_39_5_2((attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1(38
      DOWNTO 0)), attention_abs_5_qr_sva_38_0, QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_38_0,
      (RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva(38 DOWNTO 0)), attention_abs_7_qr_sva_38_0,
      STD_LOGIC_VECTOR'( RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_nor_1_ssc_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & RMS_NORM_LOOP_2_2_and_29_ssc & RMS_NORM_LOOP_2_2_and_33_ssc_1 & RMS_NORM_LOOP_2_2_and_34_ssc));
  QUANTIZE_ACTIVATION_LOOP_3_nand_seb <= NOT(CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1=STD_LOGIC_VECTOR'("11"))
      AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd);
  QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse
      <= NOT(QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1 OR QUANTIZE_ACTIVATION_LOOP_3_nand_seb);
  attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16, or_dcpl_1137);
  attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16, or_dcpl_1138);
  attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16, or_dcpl_1084);
  attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16, or_dcpl_1092);
  attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16, or_dcpl_1079);
  attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16, or_dcpl_1141);
  QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1'
      & reg_QUANTIZE_ACTIVATION_LOOP_3_quantized_value_slc_63_32_cse_slc & (APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm(55
      DOWNTO 39))) + UNSIGNED'( "00000000000000000000000001"), 26));
  QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1 <= QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_nl(25);
  attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0_mx0w6 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0, or_dcpl_1145);
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48_mx0w2 <= MUX_v_24_16_2(attention_2_1_16_16_4_4_k_proj_re_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_1_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_3_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_4_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_5_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_6_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_7_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_8_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_9_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_10_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_11_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_12_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_13_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_14_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_15_sva_1_39_16, reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2);
  attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16_mx0w5 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16, or_dcpl_1145);
  attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16, or_dcpl_1085);
  attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16, or_dcpl_1083);
  attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16, or_dcpl_1071);
  attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16, or_dcpl_1073);
  attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16, or_dcpl_1091);
  attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16, or_dcpl_1090);
  attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16, or_dcpl_1089);
  attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16, or_dcpl_1088);
  attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16, or_dcpl_1087);
  attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16, or_dcpl_1086);
  attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16, or_dcpl_1067);
  attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16, or_dcpl_1152);
  attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16, or_dcpl_1155);
  attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16, or_dcpl_1156);
  attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16, or_dcpl_1158);
  attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16, or_dcpl_1159);
  attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16, or_dcpl_1160);
  attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16, or_dcpl_1161);
  attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16, or_dcpl_1162);
  attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16, or_dcpl_1164);
  attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16, or_dcpl_1165);
  attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16, or_dcpl_1166);
  attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16, or_dcpl_1167);
  attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16, or_dcpl_1168);
  attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16, or_dcpl_1169);
  attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16, or_dcpl_1170);
  attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16, or_dcpl_1133);
  attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16, or_dcpl_1108);
  attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16, or_dcpl_1132);
  attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16, or_dcpl_1114);
  attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16, or_dcpl_1131);
  attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16, or_dcpl_1116);
  attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16, or_dcpl_1130);
  attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16, or_dcpl_1118);
  attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16, or_dcpl_1128);
  attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16, or_dcpl_1120);
  attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16, or_dcpl_1127);
  attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16, or_dcpl_1121);
  attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16, or_dcpl_1126);
  attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16, or_dcpl_1122);
  attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16, or_dcpl_1125);
  attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16, or_dcpl_1123);
  LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_7 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7, attention_2_1_16_16_4_4_quantized_hidden_states_0_6_sva_7,
      attention_2_1_16_16_4_4_quantized_hidden_states_0_7_sva_7, attention_2_1_16_16_4_4_quantized_hidden_states_0_8_sva_7,
      attention_2_1_16_16_4_4_quantized_hidden_states_0_9_sva_7, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_7, STD_LOGIC_VECTOR'( reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0));
  LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_6 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_1,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_6, STD_LOGIC_VECTOR'( reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0));
  LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_5 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_2,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_5, STD_LOGIC_VECTOR'( reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0));
  LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_4 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_3,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_4, STD_LOGIC_VECTOR'( reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0));
  LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_3 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_4,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_3, STD_LOGIC_VECTOR'( reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0));
  LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_2 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_5,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_2, STD_LOGIC_VECTOR'( reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0));
  LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_1 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_6,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_1, STD_LOGIC_VECTOR'( reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0));
  LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_0 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_7,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_0, STD_LOGIC_VECTOR'( reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0));
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_7 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7, attention_2_1_16_16_4_4_quantized_hidden_states_0_6_sva_7,
      attention_2_1_16_16_4_4_quantized_hidden_states_0_7_sva_7, attention_2_1_16_16_4_4_quantized_hidden_states_0_8_sva_7,
      attention_2_1_16_16_4_4_quantized_hidden_states_0_9_sva_7, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_7, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_6 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_1,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_6, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_5 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_2,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_5, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_4 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_3,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_4, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_3 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_4,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_3, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_2 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_5,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_2, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_1 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_6,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_1, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_0 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_7,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_0, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_7 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7, attention_2_1_16_16_4_4_quantized_hidden_states_0_6_sva_7,
      attention_2_1_16_16_4_4_quantized_hidden_states_0_7_sva_7, attention_2_1_16_16_4_4_quantized_hidden_states_0_8_sva_7,
      attention_2_1_16_16_4_4_quantized_hidden_states_0_9_sva_7, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_7, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_6 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_1,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_6, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_5 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_2,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_5, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_4 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_3,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_4, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_3 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_4,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_3, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_2 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_5,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_2, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_1 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_6,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_1, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_0 <= MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_7,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_0, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_2 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED'(
      LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1 & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0),
      2), 3) + SIGNED'( "001"), 3));
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm <= (LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_0
      AND (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_1))
      OR LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1;
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux_32_nl <= MUX_v_24_16_2(attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16, attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16, attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16, attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16, attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16, attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16, attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16, attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16, reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_7,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_7), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_1_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_6,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_6), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_3_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_1_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_2_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_5,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_5), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_4_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_2_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_3_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_4,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_4), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_5_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_3_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_4_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_3,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_3), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_6_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_4_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_5_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_2,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_2), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_7_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_5_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_6_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_1,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_1), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_8_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_6_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_7_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_0,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_0), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_9_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_7_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux_32_nl)
      + CONV_SIGNED(CONV_SIGNED(SIGNED'( LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_3_nl &
      LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_4_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_5_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_6_nl &
      LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_7_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_8_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_9_nl),
      8), 24), 24));
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1 <= LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_1
      AND (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_0);
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_1
      <= MUX_s_1_4_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7,
      STD_LOGIC_VECTOR'( reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_0
      <= MUX_s_1_4_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6,
      STD_LOGIC_VECTOR'( reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_17_nl <= MUX_v_24_16_2(attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16, attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16, attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16, attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16, attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16, attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16, attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16, attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16, reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2);
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_7,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_7), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_1_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_6,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_6), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_5_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_1_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_2_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_5,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_5), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_6_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_2_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_3_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_4,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_4), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_7_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_3_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_4_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_3,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_3), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_8_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_4_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_5_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_2,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_2), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_9_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_5_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_6_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_1,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_10_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_6_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_7_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_0,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_0), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_11_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_7_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_17_nl)
      + CONV_SIGNED(CONV_SIGNED(SIGNED'( LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_5_nl &
      LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_6_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_7_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_8_nl &
      LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_9_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_10_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_11_nl),
      8), 24), 24));
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1 <= CONV_SL_1_1(LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_conc_1_1_1_0_svs_1=STD_LOGIC_VECTOR'("10"));
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_conc_1_1_1_0_svs_1
      <= MUX_v_2_4_2((reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3(1
      DOWNTO 0)), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3(3
      DOWNTO 2)), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3(5
      DOWNTO 4)), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3(7
      DOWNTO 6)), STD_LOGIC_VECTOR'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd &
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm <= (LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_0
      AND (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_1))
      OR LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1;
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_17_nl <= MUX_v_24_16_2(attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16, attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16, attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16, attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16, attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16, attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16, attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16, attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16, reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
      & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_mux_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_7,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_7), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_mux_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_4_mux_1_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_6,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_6), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_3_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_mux_1_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_4_mux_2_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_5,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_5), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_4_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_mux_2_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_4_mux_3_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_4,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_4), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_5_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_mux_3_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_4_mux_4_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_3,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_3), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_6_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_mux_4_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_4_mux_5_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_2,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_2), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_7_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_mux_5_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_4_mux_6_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_1,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_1), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_8_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_mux_6_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  LINEAR_FORWARD_NO_MUL_LOOP_4_mux_7_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_0,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_0), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_9_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_mux_7_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_17_nl)
      + CONV_SIGNED(CONV_SIGNED(SIGNED'( LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_3_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_4_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_5_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_6_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_7_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_8_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_9_nl), 8),
      24), 24));
  LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1 <= LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_1
      AND (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_0);
  LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_1
      <= MUX_s_1_4_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7,
      STD_LOGIC_VECTOR'( LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1 & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0));
  LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_0
      <= MUX_s_1_4_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6,
      STD_LOGIC_VECTOR'( LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1 & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0));
  RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1
      <= MUX_v_24_16_2(attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16,
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_39_16, apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_3_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_re_0_7_sva_2_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_3_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_3_39_16,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1));
  GEMM_3D_FLOAT_LOOP_3_and_tmp_4_sva_mx0w2 <= GEMM_3D_FLOAT_LOOP_3_and_stg_1_3_sva_1
      AND CONV_SL_1_1(GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_0_sva_mx0w3 <= nor_1229_cse AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  GEMM_3D_FLOAT_LOOP_3_and_tmp_5_sva_mx0w2 <= GEMM_3D_FLOAT_LOOP_3_and_stg_1_2_sva_1
      AND CONV_SL_1_1(GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_1_sva_mx0w3 <= GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_1_sva_1
      AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  GEMM_3D_FLOAT_LOOP_3_and_tmp_6_sva_mx0w1 <= GEMM_3D_FLOAT_LOOP_3_and_stg_1_1_sva_1
      AND CONV_SL_1_1(GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva_mx0w3 <= GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_2_sva_1
      AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  GEMM_3D_FLOAT_LOOP_3_and_tmp_7_sva_mx0w1 <= GEMM_3D_FLOAT_LOOP_3_and_stg_1_0_sva_1
      AND CONV_SL_1_1(GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva_mx0w3 <= GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_3_sva_1
      AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1
      <= MUX_v_24_8_2(attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8
      <= MUX_v_8_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(15 DOWNTO 8)),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_8, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_15_8,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(15 DOWNTO 8)), (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(15
      DOWNTO 8)), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(15 DOWNTO 8)),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(15 DOWNTO 8)), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(15
      DOWNTO 8)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(7)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_7,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_7, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(7)),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(7)), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(7)),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(7)), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(7)),
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(6)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_6,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_6, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(6)),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(6)), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(6)),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(6)), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(6)),
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(5)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_5,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_5, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(5)),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(5)), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(5)),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(5)), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(5)),
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(4)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_4,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_4, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(4)),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(4)), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(4)),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(4)), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(4)),
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(3)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_3,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_3, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(3)),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(3)), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(3)),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(3)), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(3)),
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(2)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_2,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_2, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(2)),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(2)), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(2)),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(2)), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(2)),
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(1)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_1,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_1, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(1)),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(1)), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(1)),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(1)), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(1)),
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(0)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_0,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_0, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(0)),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(0)), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(0)),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(0)), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(0)),
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1
      <= MUX_v_24_8_2(attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_39_16, attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_39_16,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm
      <= MUX_v_8_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(15 DOWNTO 8)),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(15 DOWNTO 8)), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(7)), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(7)),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_7, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_7, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_7, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_7,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(6)), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(6)),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_6, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_6, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_6, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_6,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(5)), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(5)),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_5, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_5, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_5, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_5,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(4)), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(4)),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_4, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_4, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_4, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_4,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(3)), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(3)),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_3, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_3, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_3, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_3,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(2)), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(2)),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_2, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_2, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_2, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_2,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(1)), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(1)),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_1, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_1, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_1, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_1,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(0)), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(0)),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_0, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_0, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_0, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_0,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_1_nl
      <= MUX_v_24_8_2(attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_7_nl
      <= MUX_v_8_8_2(attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_8, reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_ftd,
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_13 & (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(12
      DOWNTO 8))), attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_8, (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0(15
      DOWNTO 8)), (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0(15 DOWNTO 8)),
      (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0(15 DOWNTO 8)), (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0(15
      DOWNTO 8)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_25_nl
      <= MUX_v_8_8_2(STD_LOGIC_VECTOR'( reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd
      & reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_1 & reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_2
      & reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_3 & reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_4
      & reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_5 & reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_6
      & reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_7), STD_LOGIC_VECTOR'(
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd & reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_1
      & reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_2 & reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_3
      & reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_4 & reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_5
      & reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_6 & reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_7),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(7 DOWNTO 0)), STD_LOGIC_VECTOR'(
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_7 & attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_6
      & attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_5 & attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_4
      & attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_3 & attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_2
      & attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_1 & attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_0),
      (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0(7 DOWNTO 0)), (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0(7
      DOWNTO 0)), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0(7 DOWNTO 0)),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0(7 DOWNTO 0)), STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED((NOT
      APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_1_nl)
      & (NOT APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_7_nl)
      & (NOT APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_25_nl))
      + SIGNED'( "0000000000000000000000000000000000000001"), 40));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_nl
      <= MUX_v_24_8_2(attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_39_16,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_6_nl
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(15)), attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_15,
      (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8(7)), (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8(7)),
      (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8(7)), (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8(7)),
      (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8(7)), (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8(7)),
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_26_nl
      <= MUX_v_3_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(14 DOWNTO 12)),
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_14_12, (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8(6
      DOWNTO 4)), (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8(6 DOWNTO 4)),
      (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8(6 DOWNTO 4)), (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8(6
      DOWNTO 4)), (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8(6 DOWNTO 4)),
      (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8(6 DOWNTO 4)), STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_27_nl
      <= MUX_v_3_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(11 DOWNTO 9)),
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_11_9, (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8(3
      DOWNTO 1)), (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8(3 DOWNTO 1)),
      (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8(3 DOWNTO 1)), (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8(3
      DOWNTO 1)), (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8(3 DOWNTO 1)),
      (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8(3 DOWNTO 1)), STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_28_nl
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(8)), attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_8,
      (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8(0)), (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8(0)),
      (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8(0)), (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8(0)),
      (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8(0)), (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8(0)),
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_16_nl
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(7)), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(7)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_7, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_7, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_7, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_7,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_17_nl
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(6)), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(6)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_6, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_6, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_6, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_6,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_18_nl
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(5)), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(5)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_5, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_5, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_5, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_5,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_19_nl
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(4)), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(4)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_4, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_4, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_4, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_4,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_20_nl
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(3)), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(3)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_3, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_3, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_3, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_3,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_21_nl
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(2)), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(2)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_2, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_2, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_2, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_2,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_22_nl
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(1)), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(1)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_1, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_1, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_1, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_1,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_23_nl
      <= MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(0)), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(0)),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_0, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_0, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_0, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_0,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED((NOT
      APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_nl)
      & (NOT APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_6_nl)
      & (NOT APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_26_nl)
      & (NOT APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_27_nl)
      & (NOT APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_28_nl)
      & (NOT APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_16_nl)
      & (NOT APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_17_nl)
      & (NOT APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_18_nl)
      & (NOT APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_19_nl)
      & (NOT APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_20_nl)
      & (NOT APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_21_nl)
      & (NOT APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_22_nl)
      & (NOT APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_23_nl))
      + SIGNED'( "0000000000000000000000000000000000000001"), 40));
  RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1
      <= MUX_v_24_16_2(attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_39_16,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1));
  RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1
      <= MUX_v_16_16_2(attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_15_0, (attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_15_8
      & attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_7 & attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_6
      & attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_5 & attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_4
      & attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_3 & attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_2
      & attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_1 & attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_0),
      attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_15_0, attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_15_0,
      attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_15_0, attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_15_0,
      attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_15_0, attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_15_0,
      attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_15_0, attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_15_0,
      (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_15_13 & attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0),
      (attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_15_8 & attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_7
      & attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_6 & attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_5
      & attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_4 & attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_3
      & attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_2 & attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_1
      & attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_0), attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_15_0,
      attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_15_0, attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_15_0,
      attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_15_0, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1));
  attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_3,
      CM_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_ctmp_sva_1, CM_LOOP_3_acc_tmp(2));
  attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx2 <= MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z(39
      DOWNTO 0)), attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_4, or_dcpl_1178);
  attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx1 <= MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z(39
      DOWNTO 0)), attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_5, or_dcpl_1180);
  attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx1 <= MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z(39
      DOWNTO 0)), attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_5, or_dcpl_1181);
  nand_378_nl <= NOT(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 AND (CM_LOOP_3_acc_tmp(0)));
  attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx1 <= MUX_v_40_2_2(CM_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_ctmp_sva_1,
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_3, nand_378_nl);
  attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx2 <= MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z(39
      DOWNTO 0)), attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_4, or_dcpl_1183);
  attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx1 <= MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z(39
      DOWNTO 0)), attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_4, or_dcpl_1184);
  attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx1 <= MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z(39
      DOWNTO 0)), attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_4, or_dcpl_1186);
  attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx1 <= MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z(39
      DOWNTO 0)), attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_4, or_dcpl_1187);
  attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_3,
      CM_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_ctmp_sva_1, CM_LOOP_3_acc_tmp(1));
  attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx2 <= MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z(39
      DOWNTO 0)), attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_4, or_dcpl_1188);
  attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx1 <= MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z(39
      DOWNTO 0)), attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_4, or_dcpl_1189);
  APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm)
      + SIGNED(APPLY_ROTARY_POS_EMB_LOOP_6_mul_3_itm), 56));
  APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1 <= APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_nl(55
      DOWNTO 16);
  APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(APPLY_ROTARY_POS_EMB_LOOP_6_mul_itm)
      + SIGNED(APPLY_ROTARY_POS_EMB_LOOP_6_mul_1_itm), 56));
  APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1 <= APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_nl(55
      DOWNTO 16);
  CACHE_UPDATE_LOOP_3_acc_sdt_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'(
      reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1),
      2), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2),
      2), 3), 3));
  TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_15_sdt_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3(2
      DOWNTO 1)), 2), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1), 2), 3), 3));
  TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_sdt_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'(
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1),
      2), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1), 2), 3), 3));
  GEMM_3D_FLOAT_LOOP_3_and_tmp_sva_mx0w0 <= GEMM_3D_FLOAT_LOOP_3_and_stg_2_3_sva_1
      AND (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2));
  GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva_mx0w0 <= GEMM_3D_FLOAT_LOOP_3_and_stg_2_0_sva_1
      AND (NOT (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2)));
  GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva_mx0w0 <= GEMM_3D_FLOAT_LOOP_3_and_stg_2_2_sva_1
      AND (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2));
  GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva_mx0w0 <= GEMM_3D_FLOAT_LOOP_3_and_stg_2_1_sva_1
      AND (NOT (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2)));
  GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva_mx0w0 <= GEMM_3D_FLOAT_LOOP_3_and_stg_2_1_sva_1
      AND (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2));
  GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva_mx0w0 <= GEMM_3D_FLOAT_LOOP_3_and_stg_2_2_sva_1
      AND (NOT (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2)));
  GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva_mx0w0 <= GEMM_3D_FLOAT_LOOP_3_and_stg_2_0_sva_1
      AND (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2));
  GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva_mx0w0 <= GEMM_3D_FLOAT_LOOP_3_and_stg_2_3_sva_1
      AND (NOT (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2)));
  GEMM_3D_FLOAT_LOOP_3_and_stg_2_0_sva_1 <= GEMM_3D_FLOAT_LOOP_3_and_stg_1_0_sva_1
      AND (NOT (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(1)));
  GEMM_3D_FLOAT_LOOP_3_and_stg_2_1_sva_1 <= GEMM_3D_FLOAT_LOOP_3_and_stg_1_1_sva_1
      AND (NOT (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(1)));
  GEMM_3D_FLOAT_LOOP_3_and_stg_2_2_sva_1 <= GEMM_3D_FLOAT_LOOP_3_and_stg_1_2_sva_1
      AND (NOT (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(1)));
  GEMM_3D_FLOAT_LOOP_3_and_stg_2_3_sva_1 <= GEMM_3D_FLOAT_LOOP_3_and_stg_1_3_sva_1
      AND (NOT (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(1)));
  GEMM_3D_FLOAT_LOOP_3_and_stg_1_0_sva_1 <= NOT((z_out_11(0)) OR (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(0)));
  GEMM_3D_FLOAT_LOOP_3_and_stg_1_1_sva_1 <= (z_out_11(0)) AND (NOT (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(0)));
  GEMM_3D_FLOAT_LOOP_3_and_stg_1_2_sva_1 <= (NOT (z_out_11(0))) AND (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(0));
  GEMM_3D_FLOAT_LOOP_3_and_stg_1_3_sva_1 <= (z_out_11(0)) AND (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(0));
  GEMM_3D_FLOAT_LOOP_4_acc_sdt_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(GEMM_3D_FLOAT_LOOP_4_acc_13_sdt_1(2
      DOWNTO 1)), 2), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1), 2), 3), 3));
  GEMM_3D_FLOAT_LOOP_4_acc_13_sdt_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(z_out_11(2
      DOWNTO 1)), 2), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1), 2), 3), 3));
  or_3014_nl <= or_dcpl_1196 OR or_dcpl_1195;
  attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6_mx1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1),40)),
      attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6, or_3014_nl);
  or_3017_nl <= or_dcpl_1199 OR or_dcpl_1198;
  attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6_mx1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1),40)),
      attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6, or_3017_nl);
  or_3019_nl <= or_dcpl_1196 OR or_dcpl_1201;
  attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6_mx1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1),40)),
      attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6, or_3019_nl);
  or_3021_nl <= or_dcpl_1199 OR or_dcpl_1203;
  attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6_mx1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1),40)),
      attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6, or_3021_nl);
  or_3022_nl <= or_dcpl_1196 OR or_dcpl_1203;
  attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6_mx1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1),40)),
      attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6, or_3022_nl);
  or_3023_nl <= or_dcpl_1199 OR or_dcpl_1201;
  attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6_mx1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1),40)),
      attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6, or_3023_nl);
  or_3024_nl <= or_dcpl_1196 OR or_dcpl_1198;
  attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6_mx1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1),40)),
      attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6, or_3024_nl);
  or_3025_nl <= or_dcpl_1199 OR or_dcpl_1195;
  attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6_mx1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1),40)),
      attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6, or_3025_nl);
  or_3027_nl <= or_dcpl_1209 OR or_dcpl_1195;
  attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6_mx1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1),40)),
      attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6, or_3027_nl);
  or_3028_nl <= or_dcpl_1209 OR or_dcpl_1198;
  attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6_mx1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1),40)),
      attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6, or_3028_nl);
  or_3029_nl <= or_dcpl_1209 OR or_dcpl_1201;
  attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6_mx1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1),40)),
      attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6, or_3029_nl);
  or_3030_nl <= or_dcpl_1209 OR or_dcpl_1203;
  attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6_mx1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1),40)),
      attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6, or_3030_nl);
  SF_LOOP_3_and_nl <= (SF_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_psp_sva_1(39))
      AND (SF_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_psp_sva_1(0));
  SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SF_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_psp_sva_1(39
      DOWNTO 1)) + CONV_SIGNED(CONV_UNSIGNED(SF_LOOP_3_and_nl, 1), 39), 39));
  SF_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_psp_sva_1 <= MUX_v_40_12_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6,
      attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6, attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6,
      attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6, attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6,
      attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6, attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6,
      attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6, attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6,
      attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6, attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6,
      attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  CM_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_ctmp_sva_1 <= MUX_v_40_4_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_3,
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_3, attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_3,
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_3, STD_LOGIC_VECTOR'( reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  CM_LOOP_3_acc_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd,
      1), 1), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1), 2), 3), 3));
  attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8_mx1 <= MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8, or_dcpl_1178);
  attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9_mx1 <= MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9, or_dcpl_1063);
  attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8_mx1 <= MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8, or_dcpl_1187);
  attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8_mx1 <= MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8, or_dcpl_1183);
  attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9_mx1 <= MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9, or_dcpl_1181);
  attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8_mx1 <= MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8, or_dcpl_1188);
  attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8_mx1 <= MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8, or_dcpl_1081);
  attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9_mx1 <= MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9, or_dcpl_1076);
  attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8_mx1 <= MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8, or_dcpl_1186);
  attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8_mx1 <= MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8, or_dcpl_1184);
  attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9_mx1 <= MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9, or_dcpl_1180);
  attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8_mx1 <= MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8, or_dcpl_1189);
  SOFTMAX_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_cse_sva_1 <= MUX_v_40_15_2(attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_3, attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_3,
      attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1,
      attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_3, attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_3,
      attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1,
      attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_3, attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_3,
      attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1,
      attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_3, attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_3,
      STD_LOGIC_VECTOR'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  operator_40_24_true_AC_TRN_AC_WRAP_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(operator_80_48_true_AC_TRN_AC_WRAP_operator_80_48_true_AC_TRN_AC_WRAP_slc_SOFTMAX_LOOP_4_sqr_56_1_itm_slc
      & (APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm(55 DOWNTO 33))) + UNSIGNED'( "000000000000000000000001"),
      24));
  SOFTMAX_LOOP_4_acc_3_cse_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(operator_40_24_true_AC_TRN_AC_WRAP_acc_nl),
      24)) & (APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm(32 DOWNTO 17))) + SIGNED(GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm),
      40));
  GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva_mx0w0 <= GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_3_sva_1
      AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva_mx0w0 <= GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_2_sva_1
      AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva_mx0w0 <= GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_1_sva_1
      AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva_mx0w0 <= nor_1229_cse AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_1_sva_1 <= reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      AND (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd);
  GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_2_sva_1 <= (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1)
      AND reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd;
  GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_3_sva_1 <= reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      AND reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd;
  GEMM_3D_FLOAT_LOOP_4_1_acc_12_sdt_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'(
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1),
      2), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2),
      2), 3), 3));
  attention_abs_5_qr_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(NOT
      (attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_2_mx0(38 DOWNTO 0))), 39),
      40) + SIGNED'( "0000000000000000000000000000000000000001"), 40));
  attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_2_mx0 <= MUX_v_40_2_2(RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1, or_dcpl_1108);
  attention_abs_6_mux_2 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(NOT
      (RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva(38 DOWNTO 0))), 39),
      40) + SIGNED'( "0000000000000000000000000000000000000001"), 40));
  QUANTIZE_ACTIVATION_LOOP_2_1_attention_abs_6_nand_nl <= NOT((attention_abs_6_mux_2(39))
      AND (RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva(39)));
  attention_abs_6_mux_3_nl <= MUX_v_39_2_2((RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva(38
      DOWNTO 0)), (attention_abs_6_mux_2(38 DOWNTO 0)), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva(39));
  QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_SIGNED(SIGNED(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      & QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_38_0), 40), 41) + CONV_UNSIGNED(CONV_SIGNED(SIGNED(QUANTIZE_ACTIVATION_LOOP_2_1_attention_abs_6_nand_nl
      & (NOT attention_abs_6_mux_3_nl)), 40), 41) + UNSIGNED'( "00000000000000000000000000000000000000001"),
      41));
  QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_itm_40_1 <= QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_nl(40);
  RMS_NORM_LOOP_2_2_and_29_ssc_1 <= (NOT QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_itm_40_1)
      AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  RMS_NORM_LOOP_2_2_and_34_ssc_1 <= (RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva(39))
      AND RMS_NORM_LOOP_2_2_and_30_m1c_1;
  RMS_NORM_LOOP_2_2_and_30_m1c_1 <= QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_itm_40_1 AND
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_nor_1_ssc_1 <= NOT((attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1(39))
      OR reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  RMS_NORM_LOOP_2_2_and_33_ssc_1 <= (NOT (RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva(39)))
      AND RMS_NORM_LOOP_2_2_and_30_m1c;
  QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1'
      & reg_QUANTIZE_ACTIVATION_LOOP_3_quantized_value_slc_63_32_cse_slc & (APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm(55
      DOWNTO 39))) + UNSIGNED'( "00000000000000000000000001"), 26));
  QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1 <= QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_nl(25);
  QUANTIZE_ACTIVATION_LOOP_3_1_nand_seb_1 <= NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      AND CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2=STD_LOGIC_VECTOR'("11"))
      AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd);
  output_0_15_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_15_lpi_4_39_16, or_dcpl_1152);
  output_0_0_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_0_lpi_4_39_16, or_dcpl_1155);
  output_0_14_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_14_lpi_4_39_16, or_dcpl_1156);
  output_0_1_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_1_lpi_4_39_16, or_dcpl_1158);
  output_0_13_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_13_lpi_4_39_16, or_dcpl_1159);
  output_0_2_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_2_lpi_4_39_16, or_dcpl_1160);
  output_0_12_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_12_lpi_4_39_16, or_dcpl_1161);
  output_0_3_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_3_lpi_4_39_16, or_dcpl_1162);
  output_0_11_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_11_lpi_4_39_16, or_dcpl_1164);
  output_0_4_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_4_lpi_4_39_16, or_dcpl_1165);
  output_0_10_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_10_lpi_4_39_16, or_dcpl_1166);
  output_0_5_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_5_lpi_4_39_16, or_dcpl_1167);
  output_0_9_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_9_lpi_4_39_16, or_dcpl_1168);
  output_0_6_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_6_lpi_4_39_16, or_dcpl_1169);
  output_0_8_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_8_lpi_4_39_16, or_dcpl_1170);
  output_0_7_lpi_4_39_16_mx1 <= MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_7_lpi_4_39_16, or_dcpl_1141);
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_7_1 <= MUX_s_1_16_2(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva,
      attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_7, attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_7,
      attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_7, attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_7,
      attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_7, attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_7,
      attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_7, attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_7,
      attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_7, attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_7,
      attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_7, attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_7,
      attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_7, attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_7,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_7, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_0_1 <= MUX_s_1_16_2(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_6_1 <= MUX_s_1_16_2(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_1_1 <= MUX_s_1_16_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_5_1 <= MUX_s_1_16_2(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_2_1 <= MUX_s_1_16_2(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_4_1 <= MUX_s_1_16_2(LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_3_1 <= MUX_s_1_16_2(reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_mux_32_nl <= MUX_v_24_16_2(output_0_0_lpi_4_39_16,
      output_0_1_lpi_4_39_16, output_0_2_lpi_4_39_16, output_0_3_lpi_4_39_16, output_0_4_lpi_4_39_16,
      output_0_5_lpi_4_39_16, output_0_6_lpi_4_39_16, output_0_7_lpi_4_39_16, output_0_8_lpi_4_39_16,
      output_0_9_lpi_4_39_16, output_0_10_lpi_4_39_16, output_0_11_lpi_4_39_16, output_0_12_lpi_4_39_16,
      output_0_13_lpi_4_39_16, output_0_14_lpi_4_39_16, output_0_15_lpi_4_39_16,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2);
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_7_1,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_7_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_1_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_6_1,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_6_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_3_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_1_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_2_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_5_1,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_5_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_4_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_2_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_3_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_4_1,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_4_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_5_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_3_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_4_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_3_1,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_3_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_6_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_4_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_5_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_2_1,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_2_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_7_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_5_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_6_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_1_1,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_1_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_8_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_6_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_7_nl <= MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_0_1,
      (NOT LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_0_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_9_nl <= LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_7_nl
      AND LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_mux_32_nl)
      + CONV_SIGNED(CONV_SIGNED(SIGNED'( LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_3_nl &
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_4_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_5_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_6_nl &
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_7_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_8_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_9_nl),
      8), 24), 24));
  CACHE_UPDATE_LOOP_2_1_acc_2_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (z_out_4(1
      DOWNTO 0))) + SIGNED'( "001"), 3));
  CACHE_UPDATE_LOOP_2_1_acc_2_itm_2_1 <= CACHE_UPDATE_LOOP_2_1_acc_2_nl(2);
  attention_max_attn_fixed_t_1_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_SIGNED(SIGNED((NOT
      reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1) & (NOT reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1)),
      40), 41) + UNSIGNED'( "00000000000000000000000000000000000000001"), 41));
  attention_max_attn_fixed_t_1_acc_1_itm_40_1 <= attention_max_attn_fixed_t_1_acc_1_nl(40);
  LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0 <= (CONV_SL_1_1(LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_conc_1_1_1_0_svs_1=STD_LOGIC_VECTOR'("01")))
      OR LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1;
  CACHE_UPDATE_LOOP_2_acc_2_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (z_out_3(1
      DOWNTO 0))) + SIGNED'( "001"), 3));
  CACHE_UPDATE_LOOP_2_acc_2_itm_2_1 <= CACHE_UPDATE_LOOP_2_acc_2_nl(2);
  SOFTMAX_LOOP_3_acc_3_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_SIGNED(SIGNED(QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39
      & QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0), 40), 41) - CONV_UNSIGNED(CONV_SIGNED(SIGNED(SOFTMAX_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_cse_sva_1),
      40), 41), 41));
  SOFTMAX_LOOP_3_acc_3_itm_40_1 <= SOFTMAX_LOOP_3_acc_3_nl(40);
  CACHE_UPDATE_LOOP_1_and_tmp <= (z_out_3(2)) AND (z_out_5(2));
  RESHAPE_2D_TO_3D_LOOP_2_2_and_cse <= (z_out_5(2)) AND (z_out_4(2));
  for_for_and_tmp <= (LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1(4)) AND LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4;
  or_dcpl_4 <= reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd OR (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  and_dcpl <= NOT((fsm_output(3)) OR (fsm_output(6)));
  and_dcpl_1 <= NOT((fsm_output(8)) OR (fsm_output(5)));
  or_tmp_11 <= (fsm_output(2)) OR (NOT (fsm_output(4)));
  nor_646_cse <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")));
  or_tmp_48 <= (NOT (fsm_output(4))) OR (fsm_output(8));
  or_dcpl_45 <= NOT((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0)) AND reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  or_dcpl_47 <= NOT(CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)=STD_LOGIC_VECTOR'("11")));
  or_dcpl_54 <= NOT(reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd AND reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  or_dcpl_60 <= (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0))) OR reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1;
  or_133_cse <= (fsm_output(4)) OR (fsm_output(8));
  or_dcpl_68 <= (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0)) OR (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  or_dcpl_79 <= (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0)) OR reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1;
  or_dcpl_96 <= (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd) OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  or_241_cse <= CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"));
  or_tmp_104 <= (fsm_output(1)) OR (fsm_output(8));
  or_255_cse <= (fsm_output(4)) OR (fsm_output(2));
  or_262_cse <= (NOT (fsm_output(1))) OR (fsm_output(8));
  mux_tmp_87 <= MUX_s_1_2_2((NOT (fsm_output(4))), (fsm_output(4)), fsm_output(2));
  mux_tmp_91 <= MUX_s_1_2_2((NOT (fsm_output(4))), (fsm_output(4)), fsm_output(5));
  nor_tmp_28 <= (fsm_output(6)) AND (fsm_output(8));
  mux_tmp_121 <= MUX_s_1_2_2((NOT (fsm_output(8))), (fsm_output(8)), fsm_output(6));
  and_dcpl_26 <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00")));
  or_349_cse <= (fsm_output(1)) OR (fsm_output(0)) OR (fsm_output(2)) OR (fsm_output(5))
      OR (fsm_output(4));
  nand_129_cse <= NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 AND
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd);
  or_361_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"));
  or_362_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_304_cse <= MUX_s_1_2_2(or_361_cse, or_362_cse, fsm_output(6));
  and_dcpl_45 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10"));
  nor_tmp_99 <= (fsm_output(4)) AND (fsm_output(8));
  and_dcpl_57 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_61 <= NOT((fsm_output(8)) OR (fsm_output(4)));
  or_619_cse <= (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd) OR (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1));
  and_dcpl_65 <= (fsm_output(1)) AND (fsm_output(3));
  or_dcpl_332 <= CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("00"));
  or_dcpl_337 <= CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("10"));
  or_dcpl_342 <= CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("01"));
  or_dcpl_351 <= NOT(CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2=STD_LOGIC_VECTOR'("11")));
  or_dcpl_377 <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd;
  or_750_cse <= (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0)) OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  or_753_cse <= (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0)) OR (NOT
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  or_tmp_330 <= NOT((fsm_output(1)) AND (fsm_output(0)) AND (fsm_output(2)) AND (NOT
      (fsm_output(4))));
  or_790_cse <= (NOT (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0)))
      OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  nand_143_cse <= NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1)));
  or_806_cse <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd OR (NOT (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1)));
  or_822_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"));
  nor_tmp_117 <= or_1984_cse AND (fsm_output(8));
  mux_tmp_363 <= MUX_s_1_2_2((fsm_output(7)), (fsm_output(8)), fsm_output(6));
  not_tmp_253 <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 4)=STD_LOGIC_VECTOR'("111")));
  or_dcpl_508 <= (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd) OR reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1;
  or_dcpl_512 <= NOT(reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd AND reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1);
  or_dcpl_584 <= reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  or_tmp_464 <= (NOT (fsm_output(6))) OR (fsm_output(8));
  nor_717_cse <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  mux_528_cse <= MUX_s_1_2_2((NOT (fsm_output(8))), (fsm_output(8)), fsm_output(4));
  or_dcpl_672 <= CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("10"));
  or_tmp_507 <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011"));
  or_1197_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100"));
  mux_tmp_604 <= MUX_s_1_2_2(or_822_cse, or_361_cse, fsm_output(6));
  mux_623_cse <= MUX_s_1_2_2((NOT (fsm_output(8))), (fsm_output(8)), fsm_output(7));
  mux_624_cse <= MUX_s_1_2_2(mux_623_cse, or_361_cse, fsm_output(6));
  or_tmp_611 <= (fsm_output(1)) OR (fsm_output(0)) OR (fsm_output(2)) OR (NOT (fsm_output(4)));
  nand_163_cse <= NOT(reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1 AND reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1);
  or_dcpl_770 <= (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2) OR
      reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0;
  or_1420_cse <= reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1 OR reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  or_dcpl_774 <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 OR reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0;
  or_1431_cse <= (NOT reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1) OR reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  or_1435_cse <= reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1 OR (NOT reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1);
  or_dcpl_791 <= NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 AND reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0);
  or_dcpl_794 <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 OR (NOT reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0);
  and_dcpl_148 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11"));
  or_tmp_682 <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("01"));
  or_dcpl_959 <= NOT((fsm_output(8)) AND (fsm_output(4)));
  or_dcpl_961 <= or_dcpl_959 OR (NOT (fsm_output(2))) OR nand_197_cse;
  and_dcpl_181 <= (NOT (fsm_output(5))) AND (fsm_output(3));
  and_dcpl_182 <= and_dcpl_181 AND and_dcpl_148;
  and_dcpl_185 <= and_dcpl_61 AND (NOT (fsm_output(2)));
  and_dcpl_186 <= and_dcpl_185 AND nor_777_cse;
  and_dcpl_187 <= and_dcpl_186 AND and_dcpl_182;
  and_dcpl_189 <= (fsm_output(5)) AND (NOT (fsm_output(3)));
  and_dcpl_190 <= and_dcpl_189 AND and_dcpl_45;
  and_dcpl_191 <= and_dcpl_61 AND (fsm_output(2));
  and_dcpl_192 <= and_dcpl_191 AND nor_777_cse;
  and_dcpl_193 <= and_dcpl_192 AND and_dcpl_190;
  and_dcpl_194 <= (fsm_output(5)) AND (fsm_output(3));
  and_dcpl_197 <= and_dcpl_186 AND and_dcpl_194 AND (NOT (z_out_5(2))) AND and_dcpl_45;
  and_dcpl_198 <= NOT((fsm_output(5)) OR (fsm_output(3)));
  and_dcpl_199 <= and_dcpl_198 AND and_dcpl_45;
  and_dcpl_200 <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_201 <= (NOT (fsm_output(8))) AND (fsm_output(4));
  and_dcpl_202 <= and_dcpl_201 AND (fsm_output(2));
  and_dcpl_203 <= and_dcpl_202 AND and_dcpl_200;
  and_dcpl_204 <= and_dcpl_203 AND and_dcpl_199;
  or_dcpl_980 <= or_dcpl_512 OR or_dcpl_4;
  or_dcpl_983 <= or_76_cse OR or_dcpl_96;
  or_dcpl_985 <= or_dcpl_508 OR or_dcpl_4;
  or_dcpl_987 <= or_130_cse OR or_dcpl_96;
  or_dcpl_988 <= or_130_cse OR or_dcpl_4;
  or_dcpl_989 <= or_dcpl_508 OR or_dcpl_96;
  or_dcpl_990 <= or_76_cse OR or_dcpl_4;
  or_dcpl_991 <= or_dcpl_512 OR or_dcpl_96;
  or_dcpl_993 <= or_dcpl_512 OR or_dcpl_584;
  or_dcpl_995 <= or_76_cse OR or_dcpl_54;
  or_dcpl_996 <= or_dcpl_508 OR or_dcpl_584;
  or_dcpl_997 <= or_130_cse OR or_dcpl_54;
  or_dcpl_998 <= or_130_cse OR or_dcpl_584;
  or_dcpl_999 <= or_dcpl_508 OR or_dcpl_54;
  or_dcpl_1000 <= or_dcpl_512 OR or_dcpl_54;
  and_dcpl_205 <= and_dcpl_201 AND (NOT (fsm_output(2)));
  and_dcpl_206 <= and_dcpl_205 AND and_dcpl_200;
  and_dcpl_207 <= and_dcpl_206 AND and_dcpl_199;
  or_dcpl_1001 <= NOT(reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 AND reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1);
  or_dcpl_1002 <= or_130_cse OR or_dcpl_1001;
  or_dcpl_1003 <= reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 OR reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  or_dcpl_1004 <= or_dcpl_508 OR or_dcpl_1003;
  or_dcpl_1005 <= (NOT reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0) OR reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  or_dcpl_1006 <= or_130_cse OR or_dcpl_1005;
  or_dcpl_1007 <= reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 OR (NOT reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1);
  or_dcpl_1008 <= or_dcpl_508 OR or_dcpl_1007;
  or_dcpl_1009 <= or_130_cse OR or_dcpl_1007;
  or_dcpl_1010 <= or_dcpl_508 OR or_dcpl_1005;
  or_dcpl_1011 <= or_130_cse OR or_dcpl_1003;
  or_dcpl_1012 <= or_dcpl_508 OR or_dcpl_1001;
  or_dcpl_1013 <= or_76_cse OR or_dcpl_1001;
  or_dcpl_1014 <= or_dcpl_512 OR or_dcpl_1003;
  or_dcpl_1015 <= or_76_cse OR or_dcpl_1005;
  or_dcpl_1016 <= or_dcpl_512 OR or_dcpl_1007;
  or_dcpl_1017 <= or_76_cse OR or_dcpl_1007;
  or_dcpl_1018 <= or_dcpl_512 OR or_dcpl_1005;
  or_dcpl_1019 <= or_dcpl_512 OR or_dcpl_1001;
  and_dcpl_209 <= and_dcpl_198 AND nor_973_cse;
  and_dcpl_211 <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_212 <= and_dcpl_205 AND and_dcpl_211;
  and_dcpl_213 <= and_dcpl_212 AND and_dcpl_199;
  nor_tmp_261 <= ((NOT((fsm_output(2)) OR (NOT (fsm_output(6))))) OR (fsm_output(4)))
      AND (fsm_output(7));
  and_dcpl_215 <= and_dcpl_202 AND and_dcpl_211;
  and_dcpl_216 <= and_dcpl_215 AND and_dcpl_199;
  mux_tmp_787 <= MUX_s_1_2_2((NOT (fsm_output(1))), (fsm_output(1)), fsm_output(0));
  mux_tmp_788 <= MUX_s_1_2_2(nand_197_cse, mux_tmp_787, fsm_output(3));
  and_dcpl_220 <= (NOT mux_tmp_788) AND and_dcpl_61 AND (NOT((fsm_output(2)) OR (fsm_output(5))))
      AND and_dcpl_148;
  and_dcpl_221 <= and_dcpl_198 AND and_dcpl_148;
  and_dcpl_222 <= and_dcpl_192 AND and_dcpl_221;
  or_dcpl_1020 <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 OR (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd);
  or_dcpl_1021 <= or_dcpl_1020 OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  or_dcpl_1022 <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd;
  or_dcpl_1023 <= or_dcpl_1022 OR (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  or_dcpl_1024 <= or_dcpl_1020 OR (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  and_dcpl_226 <= NOT((fsm_output(8)) OR (fsm_output(2)));
  or_tmp_704 <= (fsm_output(1)) OR (fsm_output(4));
  nand_253_cse <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11")));
  or_tmp_708 <= (fsm_output(3)) OR nand_253_cse;
  and_dcpl_231 <= (fsm_output(3)) AND (fsm_output(6));
  or_dcpl_1025 <= or_76_cse OR or_dcpl_584;
  and_dcpl_237 <= and_dcpl_181 AND and_dcpl_45;
  and_dcpl_239 <= and_dcpl_191 AND and_1474_cse;
  and_dcpl_240 <= and_dcpl_239 AND and_dcpl_237;
  or_dcpl_1026 <= NOT(reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd);
  or_dcpl_1027 <= (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1) OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd;
  or_dcpl_1028 <= or_dcpl_1027 OR or_dcpl_1026;
  or_dcpl_1029 <= reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 OR reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd;
  or_dcpl_1030 <= or_dcpl_1020 OR or_dcpl_1029;
  or_dcpl_1031 <= or_dcpl_1022 OR or_dcpl_1026;
  or_dcpl_1032 <= NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 AND reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd);
  or_dcpl_1033 <= or_dcpl_1032 OR or_dcpl_1029;
  or_dcpl_1034 <= (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1) OR reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd;
  or_dcpl_1035 <= or_dcpl_1027 OR or_dcpl_1034;
  or_dcpl_1036 <= reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 OR (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd);
  or_dcpl_1037 <= or_dcpl_1020 OR or_dcpl_1036;
  or_dcpl_1038 <= or_dcpl_1022 OR or_dcpl_1034;
  or_dcpl_1039 <= or_dcpl_1032 OR or_dcpl_1036;
  or_dcpl_1040 <= or_dcpl_1027 OR or_dcpl_1036;
  or_dcpl_1041 <= or_dcpl_1020 OR or_dcpl_1034;
  or_dcpl_1042 <= or_dcpl_1022 OR or_dcpl_1036;
  or_dcpl_1043 <= or_dcpl_1032 OR or_dcpl_1034;
  or_dcpl_1044 <= or_dcpl_1027 OR or_dcpl_1029;
  or_dcpl_1045 <= or_dcpl_1020 OR or_dcpl_1026;
  or_dcpl_1046 <= or_dcpl_1032 OR or_dcpl_1026;
  and_dcpl_241 <= and_dcpl_185 AND and_1474_cse;
  and_dcpl_242 <= and_dcpl_241 AND and_dcpl_209;
  and_dcpl_243 <= (fsm_output(3)) AND (NOT (fsm_output(6)));
  and_dcpl_248 <= and_dcpl_205 AND and_dcpl_200 AND (fsm_output(5)) AND and_dcpl_243
      AND (NOT (fsm_output(7))) AND (NOT((RMS_NORM_LOOP_2_2_i_4_0_sva_1(4)) AND reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1));
  and_dcpl_252 <= (fsm_output(8)) AND (NOT (fsm_output(4)));
  and_dcpl_255 <= and_dcpl_252 AND (NOT (fsm_output(2))) AND nor_777_cse AND and_dcpl_198
      AND and_dcpl_57;
  and_dcpl_256 <= and_dcpl_181 AND and_dcpl_57;
  and_dcpl_257 <= and_dcpl_239 AND and_dcpl_256;
  and_dcpl_258 <= (NOT (fsm_output(8))) AND (fsm_output(6));
  and_dcpl_259 <= and_dcpl_258 AND (NOT (fsm_output(7)));
  or_tmp_728 <= and_1559_cse OR (fsm_output(4));
  mux_817_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), or_tmp_728, fsm_output(5));
  mux_819_nl <= MUX_s_1_2_2(mux_tmp_91, mux_817_nl, fsm_output(3));
  and_dcpl_260 <= (NOT mux_819_nl) AND and_dcpl_259;
  mux_tmp_824 <= MUX_s_1_2_2(mux_tmp_121, or_2456_cse, fsm_output(4));
  nand_257_nl <= NOT((fsm_output(6)) AND (fsm_output(8)));
  mux_827_nl <= MUX_s_1_2_2(nand_257_nl, or_tmp_464, fsm_output(4));
  mux_828_nl <= MUX_s_1_2_2(mux_827_nl, or_2742_cse, fsm_output(0));
  mux_829_nl <= MUX_s_1_2_2(mux_828_nl, mux_tmp_824, fsm_output(5));
  or_1090_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"));
  mux_830_nl <= MUX_s_1_2_2(mux_829_nl, mux_2032_cse, or_1090_nl);
  mux_822_nl <= MUX_s_1_2_2(or_2742_cse, mux_2024_cse, fsm_output(0));
  mux_823_nl <= MUX_s_1_2_2(mux_822_nl, or_2736_cse, fsm_output(5));
  mux_826_nl <= MUX_s_1_2_2(mux_2032_cse, mux_823_nl, and_1773_cse);
  mux_831_nl <= MUX_s_1_2_2(mux_830_nl, mux_826_nl, fsm_output(1));
  or_dcpl_1048 <= mux_831_nl OR (fsm_output(7));
  and_dcpl_261 <= and_dcpl_181 AND nor_973_cse;
  and_dcpl_263 <= nor_tmp_99 AND (fsm_output(2));
  and_dcpl_264 <= and_dcpl_263 AND and_1474_cse;
  and_dcpl_265 <= and_dcpl_264 AND and_dcpl_261;
  or_dcpl_1050 <= NOT((fsm_output(4)) AND (fsm_output(2)));
  and_dcpl_268 <= (or_dcpl_1050 OR (NOT((fsm_output(1)) AND (fsm_output(3))))) AND
      (fsm_output(8)) AND (fsm_output(5)) AND nor_973_cse;
  and_dcpl_270 <= and_dcpl_1 AND nor_973_cse;
  mux_tmp_834 <= MUX_s_1_2_2(or_tmp_11, or_270_cse, fsm_output(1));
  mux_833_nl <= MUX_s_1_2_2(mux_tmp_87, or_270_cse, fsm_output(1));
  mux_835_nl <= MUX_s_1_2_2(mux_tmp_834, mux_833_nl, fsm_output(0));
  mux_tmp_836 <= MUX_s_1_2_2(mux_835_nl, (fsm_output(4)), fsm_output(3));
  and_dcpl_272 <= (NOT (fsm_output(8))) AND (fsm_output(2));
  and_dcpl_275 <= and_dcpl_194 AND nor_973_cse;
  and_dcpl_276 <= and_dcpl_212 AND and_dcpl_275;
  or_3137_cse <= and_1474_cse OR (fsm_output(2));
  nor_tmp_282 <= or_3137_cse AND (fsm_output(4));
  and_1498_nl <= (fsm_output(3)) AND (fsm_output(5)) AND nor_tmp_282;
  nor_897_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("000")));
  mux_837_nl <= MUX_s_1_2_2(and_1498_nl, nor_897_nl, fsm_output(6));
  and_dcpl_278 <= mux_837_nl AND and_dcpl_26;
  and_dcpl_279 <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("01"));
  or_tmp_742 <= (fsm_output(7)) OR (fsm_output(5)) OR (fsm_output(8));
  mux_tmp_839 <= MUX_s_1_2_2(or_tmp_742, or_1767_cse, fsm_output(4));
  or_1795_cse <= (fsm_output(7)) OR (NOT (fsm_output(5))) OR (fsm_output(8));
  mux_tmp_841 <= MUX_s_1_2_2(or_tmp_742, or_1795_cse, fsm_output(4));
  nor_tmp_285 <= or_3185_cse AND (fsm_output(4));
  and_dcpl_289 <= and_dcpl_202 AND nor_777_cse;
  and_dcpl_290 <= and_dcpl_289 AND and_dcpl_209;
  and_dcpl_291 <= and_dcpl_189 AND and_dcpl_148;
  and_dcpl_292 <= and_dcpl_186 AND and_dcpl_291;
  and_dcpl_293 <= and_dcpl_194 AND and_dcpl_45;
  and_dcpl_294 <= and_dcpl_239 AND and_dcpl_293;
  and_dcpl_295 <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("01"));
  or_tmp_755 <= CONV_SL_1_1(fsm_output(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("00000"));
  and_dcpl_298 <= (NOT (fsm_output(8))) AND (fsm_output(5)) AND and_dcpl_148;
  and_dcpl_302 <= and_dcpl_194 AND and_dcpl_148;
  or_tmp_757 <= nor_717_cse OR (NOT (fsm_output(4))) OR (fsm_output(8));
  or_tmp_762 <= and_1572_cse OR (fsm_output(4));
  and_337_nl <= (fsm_output(5)) AND or_tmp_762;
  mux_tmp_857 <= MUX_s_1_2_2(and_1762_cse, and_337_nl, fsm_output(3));
  mux_858_nl <= MUX_s_1_2_2(mux_tmp_857, (NOT or_tmp_755), fsm_output(6));
  and_dcpl_304 <= mux_858_nl AND and_dcpl_295;
  nor_tmp_289 <= or_1908_cse AND (fsm_output(4));
  and_dcpl_306 <= and_dcpl_264 AND and_dcpl_275;
  and_dcpl_307 <= NOT((fsm_output(8)) OR (fsm_output(6)));
  and_dcpl_308 <= and_dcpl_307 AND (NOT (fsm_output(7)));
  nor_tmp_291 <= or_1732_cse AND (fsm_output(2)) AND (fsm_output(4));
  or_tmp_767 <= and_1637_cse OR (fsm_output(4));
  and_344_nl <= (fsm_output(5)) AND or_tmp_728;
  mux_866_nl <= MUX_s_1_2_2(and_1762_cse, and_344_nl, fsm_output(3));
  nand_262_nl <= NOT((fsm_output(6)) AND mux_866_nl);
  or_1827_nl <= (fsm_output(5)) OR or_tmp_767;
  mux_865_nl <= MUX_s_1_2_2(or_2699_cse, or_1827_nl, fsm_output(3));
  or_3142_nl <= (fsm_output(6)) OR mux_865_nl;
  mux_867_nl <= MUX_s_1_2_2(nand_262_nl, or_3142_nl, fsm_output(7));
  and_dcpl_310 <= NOT(mux_867_nl OR (fsm_output(8)));
  and_dcpl_312 <= and_dcpl_185 AND and_dcpl_200;
  and_dcpl_313 <= and_dcpl_312 AND and_dcpl_190;
  and_dcpl_315 <= and_dcpl_191 AND and_dcpl_200;
  and_dcpl_316 <= and_dcpl_315 AND and_dcpl_221;
  and_dcpl_318 <= and_dcpl_202 AND and_1474_cse AND and_dcpl_199;
  and_dcpl_319 <= and_dcpl AND (fsm_output(7));
  and_dcpl_321 <= and_1474_cse AND (NOT (fsm_output(5)));
  and_dcpl_322 <= and_dcpl_202 AND and_dcpl_321;
  and_dcpl_327 <= and_dcpl_205 AND and_1474_cse;
  and_dcpl_328 <= and_dcpl_327 AND and_dcpl_237;
  or_1835_cse <= (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(5));
  and_dcpl_334 <= NOT(CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_335 <= and_dcpl_334 AND (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  and_dcpl_336 <= nor_973_cse AND (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd);
  and_dcpl_338 <= (fsm_output(0)) AND (NOT (fsm_output(5)));
  and_dcpl_339 <= and_dcpl_338 AND (NOT (fsm_output(3)));
  and_dcpl_341 <= and_dcpl_61 AND nor_717_cse;
  and_dcpl_342 <= and_dcpl_341 AND and_dcpl_339;
  nor_tmp_307 <= (fsm_output(5)) AND (fsm_output(8));
  and_dcpl_344 <= and_dcpl_206 AND and_dcpl_275;
  and_dcpl_346 <= and_dcpl_201 AND and_dcpl_211 AND and_dcpl_199;
  nand_263_cse <= NOT((fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(4)));
  or_tmp_798 <= (fsm_output(5)) OR nand_263_cse;
  mux_903_nl <= MUX_s_1_2_2(or_1867_cse, or_tmp_704, fsm_output(0));
  nand_44_nl <= NOT((fsm_output(5)) AND (NOT mux_903_nl));
  mux_904_nl <= MUX_s_1_2_2(nand_44_nl, or_tmp_798, fsm_output(3));
  and_dcpl_348 <= (NOT mux_904_nl) AND and_dcpl_272 AND and_dcpl_45;
  and_dcpl_349 <= and_dcpl_312 AND and_dcpl_293;
  and_dcpl_350 <= and_dcpl_185 AND and_dcpl_211;
  and_dcpl_351 <= and_dcpl_350 AND and_dcpl_221;
  and_dcpl_352 <= and_dcpl_241 AND and_dcpl_182;
  and_dcpl_353 <= NOT((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2)) OR (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0)));
  and_dcpl_354 <= and_dcpl_353 AND (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  and_dcpl_355 <= and_dcpl_148 AND (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(1)));
  and_dcpl_357 <= (fsm_output(0)) AND (fsm_output(5));
  and_dcpl_360 <= and_dcpl_201 AND and_1559_cse AND and_dcpl_357 AND (NOT (fsm_output(3)));
  or_dcpl_1063 <= or_dcpl_774 OR or_1420_cse;
  and_dcpl_362 <= and_dcpl_205 AND nor_777_cse;
  and_dcpl_363 <= and_dcpl_362 AND and_dcpl_275;
  and_dcpl_364 <= (fsm_output(4)) AND (NOT (fsm_output(2)));
  and_dcpl_374 <= and_dcpl_201 AND nor_717_cse AND and_dcpl_339 AND and_dcpl_45 AND
      (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1) AND (NOT(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1));
  or_tmp_805 <= (NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))))
      OR (fsm_output(8));
  mux_tmp_906 <= MUX_s_1_2_2(or_362_cse, or_361_cse, fsm_output(6));
  or_tmp_808 <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_908 <= MUX_s_1_2_2(or_1197_cse, or_tmp_808, fsm_output(4));
  mux_tmp_910 <= MUX_s_1_2_2(mux_tmp_604, or_tmp_808, fsm_output(4));
  or_tmp_812 <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_915 <= MUX_s_1_2_2(mux_tmp_906, or_tmp_812, fsm_output(4));
  or_tmp_813 <= (fsm_output(6)) OR (CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11")));
  mux_tmp_916 <= MUX_s_1_2_2(or_822_cse, (fsm_output(8)), fsm_output(6));
  mux_tmp_919 <= MUX_s_1_2_2(or_822_cse, or_362_cse, fsm_output(6));
  or_tmp_814 <= (fsm_output(6)) OR mux_623_cse;
  mux_tmp_922 <= MUX_s_1_2_2(mux_tmp_919, or_tmp_814, fsm_output(4));
  mux_tmp_927 <= MUX_s_1_2_2(mux_tmp_906, or_tmp_805, fsm_output(4));
  mux_tmp_936 <= MUX_s_1_2_2((fsm_output(7)), or_362_cse, fsm_output(6));
  mux_tmp_937 <= MUX_s_1_2_2(mux_tmp_936, or_tmp_814, fsm_output(4));
  and_dcpl_376 <= and_dcpl_191 AND and_dcpl_211;
  and_dcpl_377 <= and_dcpl_376 AND and_dcpl_293;
  or_3149_nl <= (fsm_output(6)) OR (NOT (fsm_output(2))) OR (fsm_output(4));
  or_3150_nl <= (NOT (fsm_output(6))) OR (fsm_output(2)) OR (NOT (fsm_output(4)));
  mux_953_nl <= MUX_s_1_2_2(or_3149_nl, or_3150_nl, fsm_output(7));
  and_dcpl_381 <= NOT(mux_953_nl OR (fsm_output(8)));
  and_dcpl_382 <= and_dcpl_381 AND and_dcpl_200 AND and_dcpl_198;
  or_tmp_833 <= (NOT (fsm_output(2))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  nor_923_nl <= NOT((NOT((fsm_output(2)) OR (NOT (fsm_output(4))))) OR (fsm_output(8)));
  nand_264_nl <= NOT(or_dcpl_1050 AND (fsm_output(8)));
  mux_tmp_960 <= MUX_s_1_2_2(nor_923_nl, nand_264_nl, fsm_output(1));
  mux_tmp_967 <= MUX_s_1_2_2(or_tmp_48, or_133_cse, fsm_output(2));
  or_1910_nl <= (fsm_output(2)) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_tmp_968 <= MUX_s_1_2_2(or_1910_nl, mux_tmp_967, fsm_output(1));
  and_dcpl_383 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"));
  or_1912_nl <= (fsm_output(6)) OR (NOT (fsm_output(0)));
  or_3073_nl <= (NOT (fsm_output(6))) OR (fsm_output(0));
  mux_tmp_975 <= MUX_s_1_2_2(or_1912_nl, or_3073_nl, fsm_output(7));
  and_dcpl_385 <= (NOT mux_tmp_975) AND and_dcpl_201;
  and_dcpl_386 <= and_dcpl_385 AND and_dcpl_383 AND and_dcpl_189;
  and_dcpl_388 <= and_dcpl_1 AND (fsm_output(7));
  or_tmp_861 <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(4));
  and_dcpl_390 <= and_dcpl_226 AND and_dcpl_45;
  or_tmp_878 <= NOT((fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(4)) AND (NOT
      (fsm_output(8))));
  and_dcpl_410 <= and_dcpl_376 AND and_dcpl_237;
  and_dcpl_413 <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("100"));
  nor_tmp_329 <= (fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(2)) AND (fsm_output(4));
  mux_1026_nl <= MUX_s_1_2_2((NOT nor_tmp_285), nor_tmp_329, fsm_output(5));
  mux_tmp_1027 <= MUX_s_1_2_2((NOT (fsm_output(5))), mux_1026_nl, fsm_output(3));
  and_dcpl_414 <= (NOT mux_tmp_1027) AND and_dcpl_413;
  and_dcpl_415 <= and_dcpl_312 AND and_dcpl_209;
  or_1976_nl <= (fsm_output(5)) OR (fsm_output(2)) OR (NOT (fsm_output(4)));
  or_1974_nl <= (fsm_output(5)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(2)))
      OR (fsm_output(4));
  mux_1028_nl <= MUX_s_1_2_2(or_1976_nl, or_1974_nl, fsm_output(3));
  or_tmp_913 <= (fsm_output(6)) OR mux_1028_nl;
  or_tmp_914 <= CONV_SL_1_1(fsm_output(7 DOWNTO 5)/=STD_LOGIC_VECTOR'("010"));
  and_dcpl_417 <= nor_973_cse AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd;
  and_dcpl_420 <= and_dcpl AND (NOT (fsm_output(7)));
  and_dcpl_421 <= and_dcpl_200 AND (NOT (fsm_output(5)));
  and_dcpl_422 <= and_dcpl_421 AND and_dcpl_420;
  or_dcpl_1067 <= or_619_cse OR or_750_cse;
  and_dcpl_425 <= and_dcpl_189 AND nor_973_cse;
  or_tmp_922 <= (fsm_output(4)) OR (NOT (fsm_output(7)));
  or_tmp_923 <= (NOT (fsm_output(4))) OR (fsm_output(7));
  mux_tmp_1044 <= MUX_s_1_2_2((NOT or_tmp_923), or_tmp_922, fsm_output(5));
  or_tmp_930 <= (fsm_output(5)) OR (fsm_output(4)) OR (NOT (fsm_output(7)));
  mux_tmp_1051 <= MUX_s_1_2_2(or_tmp_922, or_tmp_923, fsm_output(5));
  mux_tmp_1052 <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_923, fsm_output(5));
  or_tmp_931 <= (fsm_output(5)) OR (NOT (fsm_output(7)));
  or_dcpl_1068 <= or_dcpl_1022 OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  and_dcpl_432 <= CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1=STD_LOGIC_VECTOR'("01"));
  and_dcpl_433 <= and_dcpl_432 AND (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  or_dcpl_1070 <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd OR (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1));
  or_dcpl_1071 <= or_dcpl_1070 OR or_790_cse;
  and_dcpl_438 <= and_dcpl_203 AND and_dcpl_425;
  and_dcpl_439 <= and_dcpl_312 AND and_dcpl_256;
  or_tmp_938 <= (fsm_output(5)) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  not_tmp_549 <= NOT((fsm_output(5)) AND (fsm_output(3)) AND (fsm_output(7)));
  and_dcpl_442 <= and_dcpl_350 AND and_dcpl_293;
  and_dcpl_448 <= and_dcpl_289 AND and_dcpl_291;
  and_dcpl_449 <= nor_tmp_99 AND (NOT (fsm_output(2)));
  and_dcpl_452 <= CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1=STD_LOGIC_VECTOR'("10"));
  and_dcpl_453 <= and_dcpl_452 AND (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  or_dcpl_1073 <= nand_143_cse OR or_750_cse;
  and_dcpl_458 <= and_dcpl_353 AND reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1;
  or_dcpl_1076 <= or_dcpl_770 OR or_1435_cse;
  and_dcpl_461 <= CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1=STD_LOGIC_VECTOR'("11"));
  and_dcpl_462 <= and_dcpl_461 AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  or_dcpl_1077 <= NOT((reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0))
      AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  or_dcpl_1079 <= or_806_cse OR or_dcpl_1077;
  and_dcpl_467 <= (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2)) AND (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0));
  and_dcpl_468 <= and_dcpl_467 AND (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  or_dcpl_1081 <= or_dcpl_774 OR or_1431_cse;
  and_dcpl_471 <= and_dcpl_452 AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  or_dcpl_1083 <= nand_143_cse OR or_753_cse;
  and_dcpl_477 <= and_dcpl_385 AND nor_717_cse AND and_dcpl_194;
  and_dcpl_478 <= and_dcpl_1 AND (NOT (fsm_output(3)));
  or_tmp_992 <= nor_777_cse OR (NOT (fsm_output(2))) OR (fsm_output(4));
  mux_tmp_1113 <= MUX_s_1_2_2(or_dcpl_1050, or_tmp_11, fsm_output(1));
  or_tmp_993 <= (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(1))) OR (fsm_output(2))
      OR (fsm_output(4));
  and_dcpl_480 <= and_dcpl_334 AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  or_dcpl_1084 <= or_dcpl_1070 OR or_753_cse;
  and_dcpl_486 <= and_dcpl_461 AND (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  or_dcpl_1085 <= nand_143_cse OR or_790_cse;
  or_dcpl_1086 <= or_806_cse OR or_790_cse;
  or_dcpl_1087 <= or_619_cse OR or_753_cse;
  or_dcpl_1088 <= or_806_cse OR or_753_cse;
  or_dcpl_1089 <= or_619_cse OR or_790_cse;
  mux_tmp_1120 <= MUX_s_1_2_2(or_2456_cse, or_tmp_464, fsm_output(7));
  mux_1122_cse <= MUX_s_1_2_2(or_1197_cse, mux_tmp_1120, fsm_output(4));
  mux_1125_cse <= MUX_s_1_2_2(or_1197_cse, mux_502_cse, fsm_output(4));
  and_dcpl_511 <= (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2)) AND (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0)));
  and_dcpl_512 <= and_dcpl_511 AND (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  and_dcpl_513 <= and_dcpl_148 AND (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(1));
  or_dcpl_1090 <= or_806_cse OR or_750_cse;
  mux_1148_nl <= MUX_s_1_2_2(nand_197_cse, or_2792_cse, fsm_output(3));
  mux_1149_nl <= MUX_s_1_2_2(mux_tmp_788, mux_1148_nl, z_out_5(2));
  and_dcpl_524 <= (NOT(mux_1149_nl OR (fsm_output(8)))) AND nor_992_cse AND (NOT
      (fsm_output(5))) AND and_dcpl_148;
  nor_354_cse <= NOT((fsm_output(3)) OR (NOT (fsm_output(1))));
  nor_355_cse <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (z_out_5(2))));
  mux_1158_nl <= MUX_s_1_2_2(or_1197_cse, or_1984_cse, fsm_output(1));
  mux_1157_nl <= MUX_s_1_2_2(or_1984_cse, mux_tmp_1120, fsm_output(1));
  mux_1159_nl <= MUX_s_1_2_2(mux_1158_nl, mux_1157_nl, fsm_output(0));
  mux_1156_nl <= MUX_s_1_2_2(mux_tmp_1120, or_1197_cse, nor_355_cse);
  mux_1160_nl <= MUX_s_1_2_2(mux_1159_nl, mux_1156_nl, fsm_output(3));
  mux_1161_nl <= MUX_s_1_2_2(mux_1160_nl, mux_tmp_1120, fsm_output(2));
  mux_1154_nl <= MUX_s_1_2_2(mux_tmp_1120, mux_502_cse, nor_354_cse);
  mux_1152_nl <= MUX_s_1_2_2(mux_502_cse, mux_tmp_1120, and_1474_cse);
  mux_1153_nl <= MUX_s_1_2_2(mux_1152_nl, or_tmp_507, fsm_output(3));
  mux_1155_nl <= MUX_s_1_2_2(mux_1154_nl, mux_1153_nl, fsm_output(2));
  mux_1162_nl <= MUX_s_1_2_2(mux_1161_nl, mux_1155_nl, fsm_output(4));
  mux_tmp_1163 <= MUX_s_1_2_2(mux_1162_nl, or_tmp_507, fsm_output(5));
  and_dcpl_525 <= and_dcpl_511 AND reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1;
  and_dcpl_528 <= and_dcpl_432 AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  or_dcpl_1091 <= or_619_cse OR or_dcpl_1077;
  or_dcpl_1092 <= or_dcpl_1070 OR or_dcpl_1077;
  mux_tmp_1178 <= MUX_s_1_2_2(or_2455_cse, or_tmp_464, fsm_output(7));
  mux_tmp_1179 <= MUX_s_1_2_2(mux_tmp_1178, or_tmp_507, fsm_output(4));
  mux_tmp_1183 <= MUX_s_1_2_2((fsm_output(6)), or_tmp_464, fsm_output(7));
  mux_tmp_1185 <= MUX_s_1_2_2(or_1984_cse, mux_tmp_1183, fsm_output(4));
  mux_tmp_1187 <= MUX_s_1_2_2((fsm_output(6)), (fsm_output(8)), fsm_output(7));
  or_tmp_1035 <= and_1474_cse OR (fsm_output(3)) OR (fsm_output(8));
  and_dcpl_539 <= and_dcpl_467 AND reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1;
  or_tmp_1051 <= (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(8)));
  mux_tmp_1218 <= MUX_s_1_2_2(or_362_cse, or_822_cse, fsm_output(5));
  mux_tmp_1219 <= MUX_s_1_2_2((fsm_output(8)), or_822_cse, fsm_output(5));
  mux_tmp_1229 <= MUX_s_1_2_2(or_361_cse, or_822_cse, fsm_output(5));
  mux_tmp_1237 <= MUX_s_1_2_2(nand_253_cse, or_1984_cse, fsm_output(8));
  mux_tmp_1238 <= MUX_s_1_2_2(mux_tmp_1237, or_1197_cse, fsm_output(5));
  or_tmp_1066 <= (fsm_output(8)) OR nand_253_cse;
  mux_tmp_1240 <= MUX_s_1_2_2(or_tmp_1066, or_1197_cse, fsm_output(5));
  mux_tmp_1245 <= MUX_s_1_2_2(or_tmp_808, or_1197_cse, fsm_output(5));
  mux_1249_nl <= MUX_s_1_2_2(mux_792_cse, or_1984_cse, fsm_output(8));
  mux_tmp_1250 <= MUX_s_1_2_2(or_tmp_1066, mux_1249_nl, fsm_output(5));
  and_dcpl_548 <= and_dcpl_362 AND and_dcpl_302;
  and_dcpl_549 <= NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd OR (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(1)));
  and_dcpl_550 <= and_dcpl_549 AND (NOT (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0)));
  and_dcpl_551 <= nor_973_cse AND (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1);
  and_dcpl_552 <= and_dcpl_551 AND and_dcpl_550;
  and_dcpl_553 <= and_dcpl_338 AND (fsm_output(3));
  and_dcpl_554 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_557 <= nor_tmp_99 AND and_dcpl_554 AND and_dcpl_553 AND and_dcpl_552;
  mux_tmp_1281 <= MUX_s_1_2_2(or_255_cse, or_270_cse, fsm_output(1));
  and_dcpl_564 <= and_dcpl_198 AND (NOT (fsm_output(6)));
  and_dcpl_576 <= (fsm_output(3)) AND (NOT (fsm_output(7)));
  and_dcpl_577 <= NOT((fsm_output(1)) OR (fsm_output(5)));
  mux_1309_cse <= MUX_s_1_2_2(or_dcpl_959, or_133_cse, fsm_output(6));
  and_dcpl_581 <= and_dcpl_1 AND and_dcpl_45;
  or_tmp_1128 <= (NOT (fsm_output(1))) OR (NOT (fsm_output(2))) OR (fsm_output(4));
  and_dcpl_583 <= and_dcpl_327 AND and_dcpl_199;
  or_2235_nl <= (fsm_output(5)) OR or_tmp_762;
  mux_1311_nl <= MUX_s_1_2_2(or_2699_cse, or_2235_nl, fsm_output(3));
  or_tmp_1132 <= (fsm_output(6)) OR mux_1311_nl;
  and_443_nl <= (fsm_output(5)) AND nor_tmp_291;
  mux_1312_nl <= MUX_s_1_2_2(and_443_nl, and_1762_cse, fsm_output(3));
  nor_930_nl <= NOT((fsm_output(6)) OR mux_1312_nl);
  mux_1313_nl <= MUX_s_1_2_2(nor_930_nl, or_tmp_1132, fsm_output(7));
  or_dcpl_1104 <= mux_1313_nl OR (fsm_output(8));
  and_dcpl_585 <= and_dcpl_57 AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd;
  and_dcpl_586 <= and_dcpl_585 AND and_dcpl_486;
  and_dcpl_587 <= and_dcpl_61 AND and_dcpl_554;
  and_dcpl_588 <= and_dcpl_587 AND and_dcpl_553;
  and_dcpl_591 <= and_dcpl_57 AND (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd);
  and_dcpl_592 <= and_dcpl_591 AND and_dcpl_480;
  and_dcpl_595 <= and_dcpl_585 AND and_dcpl_471;
  and_dcpl_598 <= and_dcpl_591 AND and_dcpl_433;
  and_dcpl_601 <= and_dcpl_585 AND and_dcpl_453;
  and_dcpl_604 <= and_dcpl_591 AND and_dcpl_528;
  and_dcpl_607 <= and_dcpl_585 AND and_dcpl_528;
  and_dcpl_610 <= and_dcpl_591 AND and_dcpl_453;
  and_dcpl_613 <= and_dcpl_585 AND and_dcpl_433;
  and_dcpl_616 <= and_dcpl_591 AND and_dcpl_471;
  mux_1396_nl <= MUX_s_1_2_2(or_2249_cse, or_1983_cse, fsm_output(2));
  and_1616_nl <= (fsm_output(3)) AND (fsm_output(0)) AND (fsm_output(1));
  mux_1398_nl <= MUX_s_1_2_2(mux_806_cse, mux_1396_nl, and_1616_nl);
  mux_1399_nl <= MUX_s_1_2_2(mux_1398_nl, or_1983_cse, fsm_output(5));
  or_2296_nl <= (NOT(and_1637_cse OR (fsm_output(6)))) OR (fsm_output(7));
  mux_1394_nl <= MUX_s_1_2_2(or_2296_nl, (fsm_output(7)), fsm_output(3));
  mux_1395_nl <= MUX_s_1_2_2(or_1983_cse, mux_1394_nl, fsm_output(5));
  mux_1400_nl <= MUX_s_1_2_2(mux_1399_nl, mux_1395_nl, fsm_output(4));
  and_dcpl_618 <= NOT(mux_1400_nl OR (fsm_output(8)));
  and_dcpl_619 <= and_dcpl_241 AND and_dcpl_256;
  or_tmp_1203 <= (NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(2)) OR (NOT
      (fsm_output(4)));
  mux_1405_nl <= MUX_s_1_2_2(or_tmp_1203, or_tmp_767, fsm_output(5));
  or_2309_nl <= (fsm_output(3)) OR mux_1405_nl;
  or_1049_nl <= (NOT (fsm_output(2))) OR (fsm_output(5)) OR (fsm_output(4));
  mux_1404_nl <= MUX_s_1_2_2(or_1049_nl, or_349_cse, fsm_output(3));
  mux_1406_nl <= MUX_s_1_2_2(or_2309_nl, mux_1404_nl, fsm_output(6));
  and_dcpl_620 <= (NOT mux_1406_nl) AND and_dcpl_295;
  or_2322_nl <= (fsm_output(5)) OR or_tmp_728;
  mux_tmp_1421 <= MUX_s_1_2_2(or_2699_cse, or_2322_nl, fsm_output(3));
  or_tmp_1218 <= (fsm_output(6)) OR mux_tmp_1421;
  and_1303_nl <= (fsm_output(2)) AND (fsm_output(5)) AND (fsm_output(4));
  mux_1422_nl <= MUX_s_1_2_2(and_1303_nl, and_1762_cse, fsm_output(3));
  not_tmp_650 <= NOT((fsm_output(6)) OR mux_1422_nl);
  mux_1424_nl <= MUX_s_1_2_2(not_tmp_650, or_tmp_1132, fsm_output(7));
  mux_1423_nl <= MUX_s_1_2_2(not_tmp_650, or_tmp_1218, fsm_output(7));
  mux_1425_nl <= MUX_s_1_2_2(mux_1424_nl, mux_1423_nl, reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  and_dcpl_622 <= NOT(mux_1425_nl OR (fsm_output(8)));
  and_dcpl_625 <= (NOT((fsm_output(8)) OR (fsm_output(0)) OR (fsm_output(5)))) AND
      and_dcpl_45;
  or_tmp_1221 <= (fsm_output(1)) OR (fsm_output(2)) OR (NOT (fsm_output(4)));
  mux_tmp_1426 <= MUX_s_1_2_2(or_tmp_1221, or_tmp_1128, fsm_output(3));
  or_2328_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000"));
  mux_1427_nl <= MUX_s_1_2_2(or_2328_nl, mux_tmp_1426, reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  and_dcpl_626 <= (NOT mux_1427_nl) AND and_dcpl_625;
  and_dcpl_628 <= and_dcpl_201 AND (fsm_output(5));
  mux_1435_nl <= MUX_s_1_2_2((NOT and_1559_cse), or_3185_cse, fsm_output(3));
  nor_938_nl <= NOT((fsm_output(6)) OR mux_1435_nl);
  nor_939_nl <= NOT((NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT and_1637_cse));
  mux_1436_nl <= MUX_s_1_2_2(nor_938_nl, nor_939_nl, fsm_output(7));
  and_dcpl_629 <= mux_1436_nl AND and_dcpl_628;
  mux_tmp_1440 <= MUX_s_1_2_2((NOT and_1637_cse), or_3185_cse, fsm_output(3));
  mux_1449_nl <= MUX_s_1_2_2(and_dcpl_383, and_1559_cse, fsm_output(0));
  mux_1450_nl <= MUX_s_1_2_2((NOT or_3185_cse), mux_1449_nl, fsm_output(3));
  and_dcpl_635 <= mux_1450_nl AND (NOT (fsm_output(8))) AND (NOT (fsm_output(4)))
      AND (fsm_output(5)) AND and_dcpl_45;
  and_tmp_42 <= (fsm_output(5)) AND ((NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))))
      OR (fsm_output(4)));
  mux_tmp_1451 <= MUX_s_1_2_2(or_255_cse, or_270_cse, or_1732_cse);
  and_dcpl_641 <= and_1474_cse AND (fsm_output(5));
  and_dcpl_642 <= and_dcpl_641 AND and_dcpl_420;
  or_dcpl_1108 <= or_241_cse OR or_dcpl_79;
  or_2395_cse <= (fsm_output(5)) OR (fsm_output(2)) OR (fsm_output(4));
  mux_tmp_1489 <= MUX_s_1_2_2(or_2699_cse, or_2395_cse, fsm_output(3));
  or_dcpl_1109 <= (NOT (fsm_output(5))) OR (fsm_output(3));
  or_dcpl_1114 <= or_241_cse OR or_dcpl_68;
  and_dcpl_650 <= (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2))) AND (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0));
  and_dcpl_651 <= and_dcpl_650 AND (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  or_dcpl_1116 <= or_241_cse OR or_dcpl_60;
  and_dcpl_656 <= and_dcpl_650 AND reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1;
  or_dcpl_1118 <= or_241_cse OR or_dcpl_45;
  or_dcpl_1119 <= CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01"));
  or_dcpl_1120 <= or_dcpl_1119 OR or_dcpl_79;
  or_dcpl_1121 <= or_dcpl_1119 OR or_dcpl_68;
  or_dcpl_1122 <= or_dcpl_1119 OR or_dcpl_60;
  or_dcpl_1123 <= or_dcpl_1119 OR or_dcpl_45;
  or_dcpl_1125 <= or_dcpl_672 OR or_dcpl_79;
  or_dcpl_1126 <= or_dcpl_672 OR or_dcpl_68;
  or_dcpl_1127 <= or_dcpl_672 OR or_dcpl_60;
  or_dcpl_1128 <= or_dcpl_672 OR or_dcpl_45;
  or_dcpl_1130 <= or_dcpl_47 OR or_dcpl_79;
  or_dcpl_1131 <= or_dcpl_47 OR or_dcpl_68;
  or_dcpl_1132 <= or_dcpl_47 OR or_dcpl_60;
  or_dcpl_1133 <= or_dcpl_47 OR or_dcpl_45;
  or_tmp_1291 <= CONV_SL_1_1(fsm_output(7 DOWNTO 4)/=STD_LOGIC_VECTOR'("1000"));
  or_tmp_1296 <= (fsm_output(2)) OR (NOT (fsm_output(3))) OR (fsm_output(4)) OR (NOT
      (fsm_output(7))) OR (fsm_output(6)) OR (fsm_output(8));
  and_dcpl_718 <= and_dcpl_307 AND (fsm_output(7));
  or_tmp_1316 <= (NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("01"))))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_1519 <= MUX_s_1_2_2(or_tmp_507, or_tmp_812, fsm_output(4));
  or_tmp_1320 <= (fsm_output(3)) OR (fsm_output(4)) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(6))) OR (fsm_output(8));
  and_dcpl_721 <= and_dcpl_591 AND and_dcpl_335;
  mux_137_nl <= MUX_s_1_2_2(or_2699_cse, or_349_cse, fsm_output(3));
  not_tmp_699 <= NOT((fsm_output(6)) AND mux_137_nl);
  and_dcpl_725 <= and_dcpl_315 AND and_dcpl_256;
  and_dcpl_726 <= and_dcpl_376 AND and_dcpl_256;
  or_dcpl_1134 <= (fsm_output(5)) OR (NOT (fsm_output(3)));
  or_dcpl_1137 <= nand_143_cse OR or_dcpl_1077;
  or_dcpl_1138 <= or_dcpl_1070 OR or_750_cse;
  or_dcpl_1140 <= (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1) OR
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd;
  or_dcpl_1141 <= or_dcpl_1140 OR or_dcpl_351;
  and_dcpl_727 <= (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd) AND
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(1));
  and_dcpl_728 <= and_dcpl_727 AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0));
  and_dcpl_729 <= and_dcpl_57 AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  and_dcpl_730 <= and_dcpl_729 AND and_dcpl_728;
  and_dcpl_731 <= and_dcpl_61 AND and_dcpl_383;
  and_dcpl_732 <= and_dcpl_731 AND and_dcpl_553;
  mux_tmp_1548 <= MUX_s_1_2_2(mux_tmp_121, or_tmp_464, fsm_output(5));
  mux_tmp_1549 <= MUX_s_1_2_2(or_tmp_464, mux_tmp_121, fsm_output(5));
  nand_tmp_66 <= NOT((fsm_output(5)) AND (NOT mux_tmp_121));
  and_dcpl_735 <= and_dcpl_61 AND and_1559_cse;
  and_dcpl_736 <= and_dcpl_735 AND and_dcpl_357 AND (fsm_output(3));
  and_dcpl_739 <= and_dcpl_263 AND nor_777_cse AND and_dcpl_261;
  and_dcpl_740 <= nor_973_cse AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  and_dcpl_743 <= nor_tmp_99 AND and_dcpl_383 AND and_dcpl_553;
  and_dcpl_745 <= nor_1026_cse AND (fsm_output(3));
  and_dcpl_747 <= (NOT (fsm_output(4))) AND (fsm_output(2)) AND (fsm_output(1));
  and_dcpl_748 <= and_dcpl_747 AND and_dcpl_745;
  mux_tmp_1562 <= MUX_s_1_2_2((NOT (fsm_output(6))), (fsm_output(6)), fsm_output(7));
  and_dcpl_751 <= and_dcpl_45 AND (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(1));
  and_dcpl_753 <= and_dcpl_735 AND and_dcpl_745;
  and_dcpl_754 <= and_dcpl_753 AND and_dcpl_751 AND and_dcpl_656;
  and_dcpl_758 <= and_dcpl_45 AND (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(1)));
  and_dcpl_760 <= and_dcpl_753 AND and_dcpl_758 AND and_dcpl_512;
  and_dcpl_764 <= and_dcpl_753 AND and_dcpl_751 AND and_dcpl_651;
  and_dcpl_768 <= and_dcpl_753 AND and_dcpl_758 AND and_dcpl_525;
  and_dcpl_772 <= and_dcpl_753 AND and_dcpl_751 AND and_dcpl_458;
  and_dcpl_776 <= and_dcpl_753 AND and_dcpl_758 AND and_dcpl_468;
  and_dcpl_780 <= and_dcpl_753 AND and_dcpl_751 AND and_dcpl_354;
  and_dcpl_784 <= and_dcpl_753 AND and_dcpl_758 AND and_dcpl_539;
  and_dcpl_788 <= and_dcpl_753 AND and_dcpl_751 AND and_dcpl_512;
  and_dcpl_792 <= and_dcpl_753 AND and_dcpl_751 AND and_dcpl_525;
  and_dcpl_796 <= and_dcpl_753 AND and_dcpl_758 AND and_dcpl_458;
  and_dcpl_800 <= and_dcpl_753 AND and_dcpl_751 AND and_dcpl_468;
  and_dcpl_804 <= and_dcpl_753 AND and_dcpl_758 AND and_dcpl_354;
  and_dcpl_810 <= and_dcpl_181 AND (NOT (fsm_output(6)));
  and_dcpl_812 <= and_dcpl_376 AND and_dcpl_810 AND (fsm_output(7)) AND (LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1(4));
  and_dcpl_813 <= and_dcpl_231 AND (NOT (fsm_output(7)));
  and_dcpl_814 <= and_dcpl_747 AND and_dcpl_813;
  mux_tmp_1578 <= MUX_s_1_2_2((NOT (fsm_output(0))), (fsm_output(0)), fsm_output(5));
  and_dcpl_817 <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd AND (NOT (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(1)));
  and_dcpl_818 <= and_dcpl_817 AND (NOT (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0)));
  and_dcpl_819 <= and_dcpl_57 AND (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1);
  and_dcpl_820 <= and_dcpl_819 AND and_dcpl_818;
  and_dcpl_821 <= and_dcpl_736 AND and_dcpl_820;
  or_tmp_1354 <= (fsm_output(5)) OR (fsm_output(0));
  and_dcpl_825 <= and_dcpl_727 AND (NOT (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0)));
  and_dcpl_826 <= and_dcpl_729 AND and_dcpl_825;
  and_dcpl_827 <= and_dcpl_736 AND and_dcpl_826;
  and_dcpl_830 <= and_dcpl_817 AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0));
  and_dcpl_831 <= and_dcpl_819 AND and_dcpl_830;
  and_dcpl_832 <= and_dcpl_736 AND and_dcpl_831;
  and_dcpl_835 <= and_dcpl_549 AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0));
  and_dcpl_836 <= and_dcpl_729 AND and_dcpl_835;
  and_dcpl_837 <= and_dcpl_736 AND and_dcpl_836;
  and_dcpl_840 <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(1));
  and_dcpl_841 <= and_dcpl_840 AND (NOT (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0)));
  and_dcpl_842 <= and_dcpl_819 AND and_dcpl_841;
  and_dcpl_843 <= and_dcpl_736 AND and_dcpl_842;
  or_2500_cse <= (fsm_output(1)) OR RESHAPE_2D_TO_3D_LOOP_2_2_and_cse;
  and_dcpl_847 <= and_dcpl_205 AND or_2500_cse AND nor_1026_cse AND (NOT (fsm_output(3)))
      AND and_dcpl_45;
  and_dcpl_850 <= and_dcpl_729 AND and_dcpl_550;
  and_dcpl_851 <= and_dcpl_736 AND and_dcpl_850;
  and_dcpl_854 <= and_dcpl_840 AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0));
  and_dcpl_855 <= and_dcpl_819 AND and_dcpl_854;
  and_dcpl_856 <= and_dcpl_736 AND and_dcpl_855;
  and_dcpl_859 <= and_dcpl_729 AND and_dcpl_818;
  and_dcpl_860 <= and_dcpl_736 AND and_dcpl_859;
  and_dcpl_863 <= and_dcpl_729 AND and_dcpl_830;
  and_dcpl_864 <= and_dcpl_736 AND and_dcpl_863;
  and_dcpl_867 <= and_dcpl_819 AND and_dcpl_835;
  and_dcpl_868 <= and_dcpl_736 AND and_dcpl_867;
  and_dcpl_871 <= and_dcpl_729 AND and_dcpl_841;
  and_dcpl_872 <= and_dcpl_736 AND and_dcpl_871;
  and_dcpl_875 <= and_dcpl_819 AND and_dcpl_550;
  and_dcpl_876 <= and_dcpl_736 AND and_dcpl_875;
  and_dcpl_879 <= and_dcpl_729 AND and_dcpl_854;
  and_dcpl_880 <= and_dcpl_736 AND and_dcpl_879;
  and_dcpl_885 <= (NOT (fsm_output(5))) AND (fsm_output(7));
  or_tmp_1392 <= NOT((fsm_output(3)) AND (fsm_output(0)) AND (fsm_output(1)) AND
      (NOT (fsm_output(4))));
  and_dcpl_888 <= and_dcpl_731 AND and_dcpl_256;
  and_dcpl_959 <= and_dcpl_753 AND and_dcpl_758 AND and_dcpl_656;
  nor_946_nl <= NOT((or_2792_cse AND (fsm_output(2))) OR (fsm_output(4)));
  mux_1942_nl <= MUX_s_1_2_2(nor_946_nl, or_tmp_728, fsm_output(5));
  mux_tmp_1943 <= MUX_s_1_2_2(mux_tmp_91, mux_1942_nl, fsm_output(3));
  mux_1944_nl <= MUX_s_1_2_2(nor_992_cse, or_tmp_728, fsm_output(5));
  mux_tmp_1945 <= MUX_s_1_2_2(mux_tmp_91, mux_1944_nl, fsm_output(3));
  and_dcpl_983 <= and_dcpl_376 AND and_dcpl_810 AND (fsm_output(7)) AND (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  and_dcpl_987 <= and_dcpl_819 AND and_dcpl_825;
  and_dcpl_989 <= and_dcpl_736 AND and_dcpl_987;
  and_dcpl_999 <= and_dcpl_753 AND and_dcpl_758 AND and_dcpl_651;
  and_dcpl_1000 <= and_dcpl_819 AND and_dcpl_728;
  mux_tmp_1990 <= MUX_s_1_2_2(mux_806_cse, or_1983_cse, fsm_output(5));
  mux_tmp_1993 <= MUX_s_1_2_2(or_2249_cse, or_1983_cse, fsm_output(5));
  and_dcpl_1003 <= and_dcpl_736 AND and_dcpl_1000;
  or_dcpl_1145 <= or_76_cse OR or_dcpl_1003;
  mux_tmp_2013 <= MUX_s_1_2_2(or_1985_cse, or_tmp_914, fsm_output(4));
  mux_tmp_2015 <= MUX_s_1_2_2(or_1985_cse, or_2717_cse, fsm_output(4));
  or_dcpl_1146 <= or_dcpl_1022 OR or_dcpl_1029;
  or_2744_nl <= RESHAPE_2D_TO_3D_LOOP_2_2_and_cse OR (fsm_output(1)) OR (fsm_output(2))
      OR (NOT (fsm_output(4)));
  mux_tmp_2034 <= MUX_s_1_2_2(or_2744_nl, or_tmp_1128, fsm_output(3));
  or_2746_nl <= (fsm_output(3)) OR RESHAPE_2D_TO_3D_LOOP_2_2_and_cse OR (fsm_output(1))
      OR (fsm_output(2)) OR (NOT (fsm_output(4)));
  mux_2035_nl <= MUX_s_1_2_2(or_2746_nl, mux_tmp_2034, reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  and_dcpl_1011 <= (NOT mux_2035_nl) AND and_dcpl_625;
  and_dcpl_1033 <= and_dcpl_376 AND and_dcpl_810 AND (fsm_output(7)) AND reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  and_dcpl_1034 <= and_dcpl_362 AND and_dcpl_199;
  mux_2066_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), mux_tmp_1113, fsm_output(0));
  mux_tmp_2067 <= MUX_s_1_2_2(mux_2066_nl, or_tmp_330, fsm_output(3));
  and_dcpl_1055 <= (NOT(and_1559_cse AND (fsm_output(0)))) AND and_dcpl_201 AND and_dcpl_199;
  and_dcpl_1061 <= and_dcpl_735 AND and_dcpl_553;
  or_tmp_1632 <= and_1474_cse OR (fsm_output(2)) OR (fsm_output(4));
  or_2784_nl <= (fsm_output(5)) OR or_tmp_1632;
  mux_2085_nl <= MUX_s_1_2_2(or_2699_cse, or_2784_nl, fsm_output(3));
  not_tmp_874 <= NOT((fsm_output(6)) AND mux_2085_nl);
  or_tmp_1643 <= (NOT (fsm_output(4))) OR (fsm_output(7)) OR (fsm_output(6)) OR (NOT
      (fsm_output(8)));
  or_dcpl_1152 <= nand_129_cse OR or_dcpl_351;
  or_dcpl_1155 <= or_dcpl_377 OR or_dcpl_332;
  or_dcpl_1156 <= nand_129_cse OR or_dcpl_337;
  or_dcpl_1158 <= or_dcpl_377 OR or_dcpl_342;
  or_dcpl_1159 <= nand_129_cse OR or_dcpl_342;
  or_dcpl_1160 <= or_dcpl_377 OR or_dcpl_337;
  or_dcpl_1161 <= nand_129_cse OR or_dcpl_332;
  or_dcpl_1162 <= or_dcpl_377 OR or_dcpl_351;
  or_dcpl_1163 <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 OR (NOT
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd);
  or_dcpl_1164 <= or_dcpl_1163 OR or_dcpl_351;
  or_dcpl_1165 <= or_dcpl_1140 OR or_dcpl_332;
  or_dcpl_1166 <= or_dcpl_1163 OR or_dcpl_337;
  or_dcpl_1167 <= or_dcpl_1140 OR or_dcpl_342;
  or_dcpl_1168 <= or_dcpl_1163 OR or_dcpl_342;
  or_dcpl_1169 <= or_dcpl_1140 OR or_dcpl_337;
  or_dcpl_1170 <= or_dcpl_1163 OR or_dcpl_332;
  and_dcpl_1073 <= (NOT mux_tmp_2034) AND and_dcpl_625;
  and_dcpl_1082 <= and_dcpl_211 AND (fsm_output(5)) AND and_dcpl_813;
  and_dcpl_1084 <= or_dcpl_1138 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1088 <= or_dcpl_1084 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1091 <= or_dcpl_1071 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1094 <= or_dcpl_1092 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1097 <= or_dcpl_1090 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1100 <= or_dcpl_1088 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1103 <= or_dcpl_1086 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1106 <= or_dcpl_1079 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1109 <= or_dcpl_1067 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1112 <= or_dcpl_1087 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1115 <= or_dcpl_1089 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1118 <= or_dcpl_1091 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1121 <= or_dcpl_1073 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1124 <= or_dcpl_1083 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1127 <= or_dcpl_1085 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1130 <= or_dcpl_1137 AND and_dcpl_191 AND and_dcpl_1082;
  and_dcpl_1141 <= and_dcpl_243 AND (fsm_output(7));
  and_dcpl_1145 <= and_dcpl_279 AND and_dcpl_45;
  or_2834_cse <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01"));
  nor_953_nl <= NOT(nor_777_cse OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")));
  nor_954_nl <= NOT((fsm_output(1)) OR (fsm_output(0)) OR (fsm_output(5)) OR (NOT
      (fsm_output(6))));
  mux_2111_nl <= MUX_s_1_2_2(nor_953_nl, nor_954_nl, fsm_output(3));
  or_2833_nl <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("10"));
  mux_2110_nl <= MUX_s_1_2_2(or_2834_cse, or_2833_nl, or_1732_cse);
  nor_955_nl <= NOT((fsm_output(3)) OR mux_2110_nl);
  mux_2112_nl <= MUX_s_1_2_2(mux_2111_nl, nor_955_nl, fsm_output(2));
  nor_956_nl <= NOT((fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(1)) OR (NOT
      (fsm_output(0))) OR (fsm_output(5)) OR (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1)
      OR (fsm_output(6)));
  mux_2113_nl <= MUX_s_1_2_2(mux_2112_nl, nor_956_nl, fsm_output(4));
  and_dcpl_1151 <= mux_2113_nl AND and_dcpl_295;
  and_dcpl_1152 <= and_dcpl_186 AND and_dcpl_190;
  or_tmp_1664 <= CONV_SL_1_1(fsm_output(8 DOWNTO 5)/=STD_LOGIC_VECTOR'("1001"));
  mux_2115_nl <= MUX_s_1_2_2(or_tmp_507, or_1197_cse, fsm_output(5));
  mux_tmp_2116 <= MUX_s_1_2_2(mux_2115_nl, or_tmp_1664, fsm_output(4));
  nor_957_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(6)));
  mux_2117_nl <= MUX_s_1_2_2(nor_957_nl, and_dcpl_307, fsm_output(7));
  nand_tmp_99 <= NOT((fsm_output(5)) AND mux_2117_nl);
  mux_2118_nl <= MUX_s_1_2_2(nand_tmp_99, or_tmp_1664, fsm_output(4));
  mux_tmp_2119 <= MUX_s_1_2_2(mux_2118_nl, mux_tmp_2116, fsm_output(2));
  or_tmp_1671 <= nor_646_cse OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100"));
  mux_tmp_2121 <= MUX_s_1_2_2(mux_tmp_2119, or_tmp_1671, fsm_output(3));
  and_dcpl_1154 <= and_dcpl_449 AND and_1474_cse AND and_dcpl_261;
  and_dcpl_1162 <= and_dcpl_241 AND and_dcpl_198 AND (NOT (z_out_5(2))) AND and_dcpl_148;
  or_tmp_1690 <= (NOT (fsm_output(1))) OR (NOT (fsm_output(7))) OR (fsm_output(8));
  mux_2149_nl <= MUX_s_1_2_2(or_822_cse, mux_623_cse, nor_354_cse);
  mux_2147_nl <= MUX_s_1_2_2(mux_623_cse, or_822_cse, and_1474_cse);
  nand_286_nl <= NOT((fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(7)) AND
      (NOT (fsm_output(8))));
  mux_2148_nl <= MUX_s_1_2_2(mux_2147_nl, nand_286_nl, fsm_output(3));
  mux_2150_nl <= MUX_s_1_2_2(mux_2149_nl, mux_2148_nl, fsm_output(2));
  mux_2151_nl <= MUX_s_1_2_2(or_822_cse, mux_2150_nl, fsm_output(4));
  nand_101_nl <= NOT((fsm_output(3)) AND (NOT(nor_777_cse OR CONV_SL_1_1(fsm_output(8
      DOWNTO 7)/=STD_LOGIC_VECTOR'("01")))));
  or_2868_nl <= (fsm_output(1)) OR (NOT (fsm_output(7))) OR (fsm_output(8));
  mux_2144_nl <= MUX_s_1_2_2(or_tmp_1690, or_2868_nl, fsm_output(0));
  or_2869_nl <= (fsm_output(3)) OR mux_2144_nl;
  mux_2145_nl <= MUX_s_1_2_2(nand_101_nl, or_2869_nl, fsm_output(2));
  or_2872_nl <= (fsm_output(4)) OR mux_2145_nl;
  mux_2152_nl <= MUX_s_1_2_2(mux_2151_nl, or_2872_nl, fsm_output(5));
  or_2866_nl <= nor_355_cse OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"));
  mux_2142_nl <= MUX_s_1_2_2(or_tmp_1690, or_2866_nl, fsm_output(3));
  mux_2143_nl <= MUX_s_1_2_2(mux_2142_nl, or_361_cse, or_2395_cse);
  mux_tmp_2153 <= MUX_s_1_2_2(mux_2152_nl, mux_2143_nl, fsm_output(6));
  or_dcpl_1178 <= or_dcpl_770 OR nand_163_cse;
  nor_964_cse <= NOT((fsm_output(1)) OR (fsm_output(4)));
  mux_2172_nl <= MUX_s_1_2_2(or_1197_cse, mux_tmp_604, fsm_output(4));
  mux_2171_nl <= MUX_s_1_2_2(mux_tmp_604, mux_624_cse, fsm_output(4));
  mux_2173_nl <= MUX_s_1_2_2(mux_2172_nl, mux_2171_nl, fsm_output(1));
  or_2901_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT
      (z_out_5(2))) OR (fsm_output(4));
  mux_2170_nl <= MUX_s_1_2_2(or_1197_cse, mux_tmp_604, or_2901_nl);
  mux_2174_nl <= MUX_s_1_2_2(mux_2173_nl, mux_2170_nl, fsm_output(3));
  and_1544_nl <= nand_197_cse AND (fsm_output(4));
  mux_2168_nl <= MUX_s_1_2_2(mux_tmp_604, mux_624_cse, and_1544_nl);
  mux_2164_nl <= MUX_s_1_2_2(mux_tmp_604, or_tmp_507, fsm_output(4));
  mux_2162_nl <= MUX_s_1_2_2(or_822_cse, or_361_cse, or_1879_cse);
  mux_2165_nl <= MUX_s_1_2_2(mux_2164_nl, mux_2162_nl, and_1474_cse);
  mux_2169_nl <= MUX_s_1_2_2(mux_2168_nl, mux_2165_nl, fsm_output(3));
  mux_2175_nl <= MUX_s_1_2_2(mux_2174_nl, mux_2169_nl, fsm_output(2));
  or_2897_nl <= (NOT((NOT((NOT (fsm_output(1))) OR (fsm_output(4)))) OR (fsm_output(6))))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"));
  or_2894_nl <= (NOT(nor_964_cse OR (fsm_output(6)))) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 7)/=STD_LOGIC_VECTOR'("01"));
  mux_2160_nl <= MUX_s_1_2_2(or_2897_nl, or_2894_nl, fsm_output(0));
  or_2890_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"));
  mux_2161_nl <= MUX_s_1_2_2(mux_2160_nl, or_tmp_507, or_2890_nl);
  mux_tmp_2176 <= MUX_s_1_2_2(mux_2175_nl, mux_2161_nl, fsm_output(5));
  or_dcpl_1180 <= or_dcpl_794 OR or_1435_cse;
  or_dcpl_1181 <= or_dcpl_770 OR or_1431_cse;
  or_dcpl_1183 <= or_dcpl_770 OR or_1420_cse;
  or_dcpl_1184 <= or_dcpl_794 OR or_1420_cse;
  or_dcpl_1186 <= or_dcpl_791 OR or_1435_cse;
  or_dcpl_1187 <= or_dcpl_774 OR nand_163_cse;
  or_dcpl_1188 <= or_dcpl_774 OR or_1435_cse;
  or_dcpl_1189 <= or_dcpl_791 OR or_1420_cse;
  and_dcpl_1193 <= and_dcpl_376 AND and_dcpl_190;
  and_dcpl_1194 <= and_dcpl_239 AND and_dcpl_190;
  and_dcpl_1195 <= and_dcpl_186 AND and_dcpl_293;
  or_dcpl_1195 <= NOT((z_out_11(0)) AND (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(0)));
  or_dcpl_1196 <= CONV_SL_1_1(GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("10"));
  or_dcpl_1198 <= (z_out_11(0)) OR (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(0));
  or_dcpl_1199 <= CONV_SL_1_1(GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"));
  or_dcpl_1201 <= (z_out_11(0)) OR (NOT (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(0)));
  or_dcpl_1203 <= (NOT (z_out_11(0))) OR (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(0));
  or_dcpl_1209 <= CONV_SL_1_1(GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01"));
  and_dcpl_1199 <= and_dcpl_241 AND and_dcpl_221;
  and_1546_nl <= (fsm_output(5)) AND (fsm_output(2)) AND (fsm_output(4)) AND (NOT
      (fsm_output(8)));
  nor_968_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_2251_nl <= MUX_s_1_2_2(and_1546_nl, nor_968_nl, fsm_output(3));
  nand_tmp_104 <= NOT((fsm_output(6)) AND mux_2251_nl);
  or_3055_nl <= (fsm_output(6)) OR (NOT((NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))))
      AND (fsm_output(8))));
  mux_tmp_2252 <= MUX_s_1_2_2(or_3055_nl, nand_tmp_104, fsm_output(7));
  or_1418_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"));
  mux_2253_nl <= MUX_s_1_2_2(and_dcpl_252, (fsm_output(8)), or_1418_nl);
  nand_295_nl <= NOT(nand_240_cse AND (fsm_output(8)));
  mux_2254_nl <= MUX_s_1_2_2((NOT mux_2253_nl), nand_295_nl, fsm_output(5));
  mux_2255_nl <= MUX_s_1_2_2((NOT (fsm_output(8))), mux_2254_nl, fsm_output(3));
  or_3058_nl <= (fsm_output(6)) OR mux_2255_nl;
  mux_2256_itm <= MUX_s_1_2_2(or_3058_nl, nand_tmp_104, fsm_output(7));
  and_dcpl_1225 <= and_dcpl_263 AND and_dcpl_211 AND and_dcpl_275;
  and_dcpl_1227 <= and_dcpl_263 AND and_dcpl_200 AND and_dcpl_261;
  and_1550_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"));
  nor_969_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")));
  mux_2259_nl <= MUX_s_1_2_2(and_1550_nl, nor_969_nl, fsm_output(6));
  and_dcpl_1232 <= mux_2259_nl AND CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("10"));
  mux_868_nl <= MUX_s_1_2_2(or_dcpl_1050, nor_tmp_282, fsm_output(5));
  mux_869_nl <= MUX_s_1_2_2(mux_868_nl, mux_tmp_91, fsm_output(3));
  rms_norm_16_div_cmp_a_mx0c0 <= (NOT mux_869_nl) AND and_dcpl_308;
  attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c0 <= and_dcpl_342 AND and_dcpl_336
      AND and_dcpl_335;
  attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c9 <= and_dcpl_360 AND and_dcpl_355
      AND and_dcpl_354;
  nor_998_cse <= NOT(nor_777_cse OR (fsm_output(4)));
  nor_999_nl <= NOT((NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (fsm_output(4))
      OR (fsm_output(8)));
  mux_1007_nl <= MUX_s_1_2_2(nor_999_nl, (fsm_output(8)), fsm_output(5));
  mux_1008_nl <= MUX_s_1_2_2((NOT mux_1007_nl), mux_958_cse, fsm_output(6));
  nand_322_nl <= NOT(or_1732_cse AND (fsm_output(4)) AND (fsm_output(8)));
  nor_1001_nl <= NOT(nor_176_cse OR (fsm_output(8)));
  mux_1005_nl <= MUX_s_1_2_2(nand_322_nl, nor_1001_nl, fsm_output(5));
  or_1952_nl <= nor_964_cse OR (fsm_output(8));
  or_1950_nl <= (NOT((NOT LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4) OR (NOT (fsm_output(1)))
      OR (fsm_output(4)))) OR (fsm_output(8));
  mux_1003_nl <= MUX_s_1_2_2(or_1952_nl, or_1950_nl, fsm_output(0));
  mux_1004_nl <= MUX_s_1_2_2(mux_1003_nl, or_133_cse, fsm_output(5));
  mux_1006_nl <= MUX_s_1_2_2(mux_1005_nl, mux_1004_nl, fsm_output(6));
  mux_1009_nl <= MUX_s_1_2_2(mux_1008_nl, mux_1006_nl, fsm_output(3));
  nand_323_nl <= NOT((fsm_output(5)) AND ((or_1732_cse AND (fsm_output(4))) OR (fsm_output(8))));
  mux_1001_nl <= MUX_s_1_2_2(nand_323_nl, mux_958_cse, fsm_output(6));
  nand_325_nl <= NOT(nand_263_cse AND (fsm_output(8)));
  mux_998_nl <= MUX_s_1_2_2(or_dcpl_959, nand_325_nl, fsm_output(5));
  or_1944_nl <= (fsm_output(1)) OR (fsm_output(4)) OR (fsm_output(8));
  mux_997_nl <= MUX_s_1_2_2((fsm_output(8)), or_1944_nl, fsm_output(5));
  mux_999_nl <= MUX_s_1_2_2(mux_998_nl, mux_997_nl, fsm_output(6));
  mux_1002_nl <= MUX_s_1_2_2(mux_1001_nl, mux_999_nl, fsm_output(3));
  mux_1010_nl <= MUX_s_1_2_2(mux_1009_nl, mux_1002_nl, fsm_output(2));
  mux_993_nl <= MUX_s_1_2_2(or_tmp_878, (fsm_output(8)), fsm_output(5));
  or_1943_nl <= (fsm_output(5)) OR (fsm_output(1)) OR (fsm_output(4)) OR (fsm_output(8));
  mux_994_nl <= MUX_s_1_2_2(mux_993_nl, or_1943_nl, fsm_output(6));
  mux_991_nl <= MUX_s_1_2_2(or_tmp_878, or_tmp_48, fsm_output(5));
  or_1940_nl <= (NOT (fsm_output(5))) OR (fsm_output(0)) OR (fsm_output(1)) OR (NOT
      (fsm_output(4))) OR (fsm_output(8));
  mux_992_nl <= MUX_s_1_2_2(mux_991_nl, or_1940_nl, fsm_output(6));
  mux_995_nl <= MUX_s_1_2_2(mux_994_nl, mux_992_nl, fsm_output(3));
  or_1939_nl <= (fsm_output(1)) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  or_1938_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_987_nl <= MUX_s_1_2_2(or_1939_nl, or_1938_nl, fsm_output(0));
  or_1937_nl <= nor_998_cse OR (fsm_output(8));
  mux_988_nl <= MUX_s_1_2_2(mux_987_nl, or_1937_nl, fsm_output(5));
  or_1934_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_989_nl <= MUX_s_1_2_2(mux_988_nl, or_1934_nl, fsm_output(6));
  or_1932_nl <= (fsm_output(0)) OR (NOT (fsm_output(1))) OR (fsm_output(4)) OR (fsm_output(8));
  or_1931_nl <= (NOT((fsm_output(0)) OR (NOT (fsm_output(1))) OR (fsm_output(4))))
      OR (fsm_output(8));
  mux_986_nl <= MUX_s_1_2_2(or_1932_nl, or_1931_nl, fsm_output(5));
  or_1933_nl <= (fsm_output(6)) OR mux_986_nl;
  mux_990_nl <= MUX_s_1_2_2(mux_989_nl, or_1933_nl, fsm_output(3));
  mux_996_nl <= MUX_s_1_2_2(mux_995_nl, mux_990_nl, fsm_output(2));
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c0 <= MUX_s_1_2_2(mux_1010_nl,
      mux_996_nl, fsm_output(7));
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c2 <= (NOT((CONV_SL_1_1(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0=STD_LOGIC_VECTOR'("1111"))
      AND LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4) OR mux_tmp_975)) AND and_dcpl_202
      AND (NOT (fsm_output(1))) AND (fsm_output(5)) AND (NOT (fsm_output(3)));
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c3 <= (NOT(mux_tmp_975 OR (fsm_output(8))))
      AND and_1771_cse AND (NOT (fsm_output(1))) AND and_dcpl_189 AND LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4
      AND CONV_SL_1_1(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0=STD_LOGIC_VECTOR'("1111"));
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c5 <= and_dcpl_241 AND and_dcpl_181
      AND (fsm_output(6)) AND (NOT((fsm_output(7)) OR LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4));
  mux_1022_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), (fsm_output(6)), fsm_output(5));
  mux_1023_nl <= MUX_s_1_2_2(mux_1022_nl, or_2834_cse, fsm_output(1));
  nor_1019_nl <= NOT((fsm_output(3)) OR mux_1023_nl);
  nor_1020_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(5))) OR (fsm_output(6)));
  nor_1021_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(5))) OR (fsm_output(6)));
  mux_1021_nl <= MUX_s_1_2_2(nor_1020_nl, nor_1021_nl, fsm_output(0));
  mux_1024_nl <= MUX_s_1_2_2(nor_1019_nl, mux_1021_nl, fsm_output(2));
  nor_1022_nl <= NOT((NOT(and_1474_cse OR (fsm_output(5)))) OR (fsm_output(6)));
  nor_1023_nl <= NOT((NOT((NOT((fsm_output(3)) OR (fsm_output(1)))) OR (fsm_output(5))))
      OR (fsm_output(6)));
  nor_1024_nl <= NOT((NOT(nor_354_cse OR (fsm_output(5)))) OR (fsm_output(6)));
  mux_1019_nl <= MUX_s_1_2_2(nor_1023_nl, nor_1024_nl, fsm_output(0));
  mux_1020_nl <= MUX_s_1_2_2(nor_1022_nl, mux_1019_nl, fsm_output(2));
  mux_1025_nl <= MUX_s_1_2_2(mux_1024_nl, mux_1020_nl, fsm_output(4));
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c7 <= mux_1025_nl AND and_dcpl_295;
  mux_1029_nl <= MUX_s_1_2_2(or_tmp_728, or_tmp_704, fsm_output(0));
  mux_1030_nl <= MUX_s_1_2_2((NOT mux_1029_nl), or_tmp_767, fsm_output(5));
  mux_1031_nl <= MUX_s_1_2_2(mux_tmp_91, mux_1030_nl, fsm_output(3));
  nand_49_nl <= NOT((fsm_output(6)) AND (NOT mux_1031_nl));
  mux_1032_nl <= MUX_s_1_2_2(nand_49_nl, or_tmp_913, fsm_output(7));
  for_for_strm_in_tmp_sva_31_2_mx0c1 <= NOT(mux_1032_nl OR (fsm_output(8)));
  GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c0 <= and_dcpl_342 AND and_dcpl_417 AND and_dcpl_335;
  GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c1 <= or_dcpl_1067 AND and_dcpl_185 AND and_dcpl_422;
  GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c2 <= and_dcpl_289 AND and_dcpl_425;
  GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c4 <= and_dcpl_186 AND and_dcpl_256;
  GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c7 <= and_dcpl_192 AND and_dcpl_293;
  GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c9 <= and_dcpl_315 AND and_dcpl_182;
  GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c10 <= and_dcpl_327 AND and_dcpl_291;
  attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c0 <= and_dcpl_342 AND and_dcpl_417
      AND and_dcpl_453;
  attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c1 <= or_dcpl_1073 AND and_dcpl_185
      AND and_dcpl_422;
  nor_1031_nl <= NOT((NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))))
      OR (fsm_output(8)));
  nand_330_nl <= NOT((NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"))))
      AND (fsm_output(8)));
  mux_1078_nl <= MUX_s_1_2_2(nor_1031_nl, nand_330_nl, fsm_output(4));
  or_2029_cse <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00")) OR
      mux_1078_nl;
  or_3163_cse <= (z_out_5(2)) OR (fsm_output(0));
  nor_1032_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(1)))
      OR (fsm_output(8)));
  nor_1033_nl <= NOT((fsm_output(3)) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(8)));
  mux_1076_nl <= MUX_s_1_2_2(nor_1032_nl, nor_1033_nl, fsm_output(2));
  nand_50_cse <= NOT((NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("01"))))
      AND mux_1076_nl);
  or_2022_nl <= (or_3163_cse AND (fsm_output(1))) OR (fsm_output(8));
  mux_1073_nl <= MUX_s_1_2_2(or_1848_cse, or_2022_nl, fsm_output(3));
  mux_1074_cse <= MUX_s_1_2_2(mux_1073_nl, (fsm_output(8)), or_255_cse);
  or_2019_nl <= (NOT(CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)/=STD_LOGIC_VECTOR'("00")) OR (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1)
      OR (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0)) OR CONV_SL_1_1(fsm_output(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10111")))) OR (fsm_output(8));
  mux_1075_nl <= MUX_s_1_2_2(mux_1074_cse, or_2019_nl, fsm_output(5));
  mux_1077_nl <= MUX_s_1_2_2(nand_50_cse, mux_1075_nl, fsm_output(6));
  mux_1079_itm <= MUX_s_1_2_2(or_2029_cse, mux_1077_nl, fsm_output(7));
  mux_1088_nl <= MUX_s_1_2_2(or_tmp_104, or_262_cse, fsm_output(0));
  mux_1089_cse <= MUX_s_1_2_2(mux_1088_nl, (fsm_output(8)), or_2797_cse);
  or_2038_nl <= nor_355_cse OR (fsm_output(8));
  mux_1085_nl <= MUX_s_1_2_2(or_262_cse, or_2038_nl, fsm_output(3));
  mux_1086_nl <= MUX_s_1_2_2(mux_1085_nl, (fsm_output(8)), fsm_output(4));
  nand_52_nl <= NOT((fsm_output(7)) AND (NOT mux_1086_nl));
  mux_1087_cse <= MUX_s_1_2_2(nand_52_nl, or_361_cse, fsm_output(5));
  nand_332_nl <= NOT(nand_381_cse AND (fsm_output(8)));
  nor_1035_nl <= NOT(and_1474_cse OR (fsm_output(8)));
  nor_1036_nl <= NOT((NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (fsm_output(8)));
  mux_1081_nl <= MUX_s_1_2_2(nor_1035_nl, nor_1036_nl, fsm_output(3));
  nand_51_nl <= NOT((fsm_output(4)) AND mux_1081_nl);
  mux_1082_nl <= MUX_s_1_2_2(nand_332_nl, nand_51_nl, fsm_output(7));
  mux_1080_nl <= MUX_s_1_2_2(or_262_cse, or_tmp_104, fsm_output(0));
  or_2034_nl <= (NOT (fsm_output(7))) OR (fsm_output(4)) OR (fsm_output(3)) OR mux_1080_nl;
  mux_1083_nl <= MUX_s_1_2_2(mux_1082_nl, or_2034_nl, fsm_output(5));
  mux_1084_cse <= MUX_s_1_2_2(mux_1083_nl, or_361_cse, fsm_output(6));
  or_2039_nl <= (NOT (fsm_output(4))) OR (fsm_output(3)) OR (NOT (fsm_output(0)))
      OR (NOT (fsm_output(1))) OR (fsm_output(8));
  mux_1090_nl <= MUX_s_1_2_2((NOT mux_1089_cse), or_2039_nl, fsm_output(7));
  or_2041_nl <= (fsm_output(5)) OR mux_1090_nl;
  mux_1091_nl <= MUX_s_1_2_2(or_2041_nl, mux_1087_cse, fsm_output(6));
  attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c7 <= MUX_s_1_2_2(mux_1091_nl,
      mux_1084_cse, fsm_output(2));
  attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c9 <= and_dcpl_360 AND and_dcpl_355
      AND and_dcpl_458;
  attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c0 <= and_dcpl_342 AND and_dcpl_336
      AND and_dcpl_462;
  attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c1 <= or_dcpl_1079 AND and_dcpl_185
      AND and_dcpl_422;
  or_2068_nl <= (NOT (fsm_output(4))) OR (fsm_output(3)) OR (NOT (fsm_output(1)))
      OR (fsm_output(8));
  mux_1110_nl <= MUX_s_1_2_2((NOT mux_1089_cse), or_2068_nl, fsm_output(7));
  or_2070_nl <= (fsm_output(5)) OR mux_1110_nl;
  mux_1111_nl <= MUX_s_1_2_2(or_2070_nl, mux_1087_cse, fsm_output(6));
  attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c7 <= MUX_s_1_2_2(mux_1111_nl,
      mux_1084_cse, fsm_output(2));
  attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c9 <= and_dcpl_360 AND and_dcpl_355
      AND and_dcpl_468;
  apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c0 <= and_dcpl_342 AND and_dcpl_417
      AND and_dcpl_471;
  apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c1 <= or_dcpl_1083 AND and_dcpl_185
      AND and_dcpl_422;
  attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c0 <= and_dcpl_342 AND and_dcpl_417
      AND and_dcpl_433;
  attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c1 <= or_dcpl_1089 AND and_dcpl_185
      AND and_dcpl_422;
  mux_1129_nl <= MUX_s_1_2_2(mux_1125_cse, mux_tmp_1120, fsm_output(0));
  mux_1130_nl <= MUX_s_1_2_2(mux_1122_cse, mux_1129_nl, fsm_output(2));
  mux_1126_nl <= MUX_s_1_2_2(or_1984_cse, mux_tmp_1120, fsm_output(4));
  mux_1127_nl <= MUX_s_1_2_2(mux_1126_nl, mux_1125_cse, fsm_output(0));
  mux_1128_nl <= MUX_s_1_2_2(mux_1127_nl, mux_tmp_1120, fsm_output(2));
  mux_1131_nl <= MUX_s_1_2_2(mux_1130_nl, mux_1128_nl, fsm_output(1));
  mux_1121_nl <= MUX_s_1_2_2(mux_tmp_1120, or_tmp_507, fsm_output(4));
  mux_1123_nl <= MUX_s_1_2_2(mux_1122_cse, mux_1121_nl, fsm_output(2));
  mux_1132_cse <= MUX_s_1_2_2(mux_1131_nl, mux_1123_nl, fsm_output(3));
  attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c5 <= and_dcpl_185 AND ((fsm_output(1))
      XOR (fsm_output(3))) AND and_dcpl_338 AND and_dcpl_148;
  attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c8 <= and_dcpl_350 AND and_dcpl_182;
  attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c10 <= and_dcpl_360 AND and_dcpl_513
      AND and_dcpl_512;
  attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c0 <= and_dcpl_342 AND and_dcpl_336
      AND and_dcpl_453;
  attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c1 <= or_dcpl_1090 AND and_dcpl_185
      AND and_dcpl_422;
  or_2095_nl <= (CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
      AND reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 AND (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0)))
      AND CONV_SL_1_1(fsm_output(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"))) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("011"));
  mux_1147_itm <= MUX_s_1_2_2(mux_1132_cse, or_2095_nl, fsm_output(5));
  attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c10 <= and_dcpl_360 AND and_dcpl_513
      AND and_dcpl_525;
  attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c0 <= and_dcpl_342 AND and_dcpl_417
      AND and_dcpl_528;
  attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c1 <= or_dcpl_1091 AND and_dcpl_185
      AND and_dcpl_422;
  or_2110_nl <= (CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
      AND (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) AND (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0))
      AND CONV_SL_1_1(fsm_output(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"))) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("011"));
  mux_1177_itm <= MUX_s_1_2_2(mux_1132_cse, or_2110_nl, fsm_output(5));
  attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c10 <= and_dcpl_360 AND and_dcpl_513
      AND and_dcpl_468;
  attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c0 <= and_dcpl_342 AND and_dcpl_336
      AND and_dcpl_528;
  attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c1 <= or_dcpl_1092 AND and_dcpl_185
      AND and_dcpl_422;
  mux_1193_nl <= MUX_s_1_2_2(or_1197_cse, mux_tmp_1183, fsm_output(4));
  mux_1191_nl <= MUX_s_1_2_2(or_1984_cse, mux_tmp_1187, fsm_output(4));
  mux_1192_nl <= MUX_s_1_2_2(mux_1191_nl, mux_tmp_1183, fsm_output(0));
  mux_1194_nl <= MUX_s_1_2_2(mux_1193_nl, mux_1192_nl, fsm_output(2));
  mux_1188_nl <= MUX_s_1_2_2(or_1197_cse, mux_tmp_1187, fsm_output(4));
  mux_1189_nl <= MUX_s_1_2_2(mux_tmp_1185, mux_1188_nl, fsm_output(0));
  mux_1190_nl <= MUX_s_1_2_2(mux_1189_nl, mux_tmp_1183, fsm_output(2));
  mux_1195_nl <= MUX_s_1_2_2(mux_1194_nl, mux_1190_nl, fsm_output(1));
  mux_1184_nl <= MUX_s_1_2_2(mux_tmp_1183, mux_tmp_1178, fsm_output(4));
  mux_1186_nl <= MUX_s_1_2_2(mux_tmp_1185, mux_1184_nl, fsm_output(2));
  mux_1196_nl <= MUX_s_1_2_2(mux_1195_nl, mux_1186_nl, fsm_output(3));
  or_2121_nl <= (fsm_output(4)) OR mux_tmp_1178;
  and_1593_nl <= CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
      AND reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 AND (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0));
  mux_1180_nl <= MUX_s_1_2_2(mux_tmp_1179, or_2121_nl, and_1593_nl);
  mux_1181_nl <= MUX_s_1_2_2(mux_tmp_1178, mux_1180_nl, and_1572_cse);
  mux_1182_nl <= MUX_s_1_2_2(mux_1181_nl, mux_tmp_1179, fsm_output(3));
  mux_1197_itm <= MUX_s_1_2_2(mux_1196_nl, mux_1182_nl, fsm_output(5));
  nor_1043_nl <= NOT((fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(0)) OR (fsm_output(3))
      OR (fsm_output(8)));
  and_1595_nl <= (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(8));
  mux_1205_nl <= MUX_s_1_2_2(nor_1043_nl, and_1595_nl, fsm_output(4));
  or_2130_nl <= (or_2792_cse AND (fsm_output(3))) OR (fsm_output(8));
  mux_1203_nl <= MUX_s_1_2_2(or_2130_nl, or_tmp_1035, fsm_output(2));
  mux_1204_nl <= MUX_s_1_2_2((fsm_output(8)), mux_1203_nl, fsm_output(4));
  mux_1206_nl <= MUX_s_1_2_2(mux_1205_nl, mux_1204_nl, fsm_output(5));
  or_2132_nl <= (fsm_output(6)) OR mux_1206_nl;
  or_2129_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(8));
  mux_1201_nl <= MUX_s_1_2_2(or_2129_nl, or_tmp_1035, fsm_output(2));
  or_3166_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("01")) OR mux_1201_nl;
  or_2127_nl <= (NOT (fsm_output(3))) OR (fsm_output(8));
  or_2126_nl <= (z_out_5(2)) OR (NOT (fsm_output(3))) OR (fsm_output(8));
  mux_1198_nl <= MUX_s_1_2_2(or_2126_nl, (fsm_output(8)), fsm_output(0));
  mux_1199_nl <= MUX_s_1_2_2(or_2127_nl, mux_1198_nl, fsm_output(1));
  mux_1200_nl <= MUX_s_1_2_2(mux_1199_nl, (fsm_output(8)), or_2395_cse);
  mux_1202_nl <= MUX_s_1_2_2(or_3166_nl, mux_1200_nl, fsm_output(6));
  attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c10 <= MUX_s_1_2_2(or_2132_nl,
      mux_1202_nl, fsm_output(7));
  attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c12 <= and_dcpl_360 AND and_dcpl_513
      AND and_dcpl_539;
  or_2184_nl <= and_1771_cse OR (fsm_output(8));
  mux_1270_nl <= MUX_s_1_2_2(mux_tmp_967, or_2184_nl, fsm_output(1));
  mux_1271_nl <= MUX_s_1_2_2(mux_tmp_968, mux_1270_nl, fsm_output(0));
  nor_1050_nl <= NOT(nor_tmp_291 OR (fsm_output(8)));
  mux_1272_nl <= MUX_s_1_2_2(mux_1271_nl, nor_1050_nl, fsm_output(5));
  mux_1268_nl <= MUX_s_1_2_2(and_dcpl_61, mux_528_cse, or_3185_cse);
  mux_1267_nl <= MUX_s_1_2_2((NOT (fsm_output(8))), mux_tmp_960, fsm_output(0));
  mux_1269_nl <= MUX_s_1_2_2((NOT mux_1268_nl), mux_1267_nl, fsm_output(5));
  mux_1273_nl <= MUX_s_1_2_2(mux_1272_nl, mux_1269_nl, fsm_output(3));
  nor_1325_nl <= NOT((fsm_output(6)) OR mux_1273_nl);
  nor_1326_nl <= NOT((fsm_output(5)) OR and_1474_cse OR (fsm_output(2)) OR (NOT (fsm_output(4)))
      OR (fsm_output(8)));
  nor_1327_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(1))) OR (fsm_output(2))
      OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1265_nl <= MUX_s_1_2_2(nor_1326_nl, nor_1327_nl, fsm_output(3));
  nor_1328_nl <= NOT(nor_1106_cse OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  nor_1329_nl <= NOT(and_1474_cse OR (NOT (fsm_output(2))) OR (NOT (fsm_output(4)))
      OR (fsm_output(8)));
  mux_1263_nl <= MUX_s_1_2_2(nor_1328_nl, nor_1329_nl, fsm_output(5));
  nor_1330_nl <= NOT((NOT(and_1572_cse OR (fsm_output(4)))) OR (fsm_output(8)));
  nor_1331_nl <= NOT((fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(2)) OR (NOT
      (fsm_output(4))) OR (fsm_output(8)));
  mux_1262_nl <= MUX_s_1_2_2(nor_1330_nl, nor_1331_nl, fsm_output(5));
  mux_1264_nl <= MUX_s_1_2_2(mux_1263_nl, mux_1262_nl, fsm_output(3));
  mux_1266_nl <= MUX_s_1_2_2(mux_1265_nl, mux_1264_nl, fsm_output(6));
  GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c0 <= MUX_s_1_2_2(nor_1325_nl, mux_1266_nl,
      fsm_output(7));
  nor_1053_cse <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (fsm_output(1))
      OR (NOT (fsm_output(2))) OR (fsm_output(4)));
  nor_1054_nl <= NOT((fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(1)))
      OR (fsm_output(2)) OR (NOT (fsm_output(4))));
  mux_1275_nl <= MUX_s_1_2_2(nor_1053_cse, nor_1054_nl, fsm_output(7));
  nor_1055_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0)))
      OR (fsm_output(1)) OR (NOT (fsm_output(2))) OR (fsm_output(4)));
  mux_1276_nl <= MUX_s_1_2_2(mux_1275_nl, nor_1055_nl, CACHE_UPDATE_LOOP_1_and_tmp);
  GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c1 <= mux_1276_nl AND and_dcpl_1 AND (fsm_output(3));
  or_2199_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(2))) OR (fsm_output(0))
      OR (NOT (fsm_output(6))) OR (fsm_output(7));
  or_2198_nl <= (fsm_output(2)) OR (fsm_output(0)) OR (fsm_output(6)) OR (NOT (fsm_output(7)));
  mux_1279_nl <= MUX_s_1_2_2(or_2199_nl, or_2198_nl, fsm_output(5));
  or_3169_nl <= (fsm_output(4)) OR mux_1279_nl;
  or_2195_nl <= (NOT (fsm_output(2))) OR (fsm_output(0)) OR (fsm_output(6)) OR (NOT
      (fsm_output(7)));
  or_2193_nl <= (NOT CACHE_UPDATE_LOOP_1_and_tmp) OR (fsm_output(0)) OR (fsm_output(6))
      OR (NOT (fsm_output(7)));
  mux_1277_nl <= MUX_s_1_2_2(or_2193_nl, or_2249_cse, fsm_output(2));
  mux_1278_nl <= MUX_s_1_2_2(or_2195_nl, mux_1277_nl, fsm_output(3));
  or_3170_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("01")) OR mux_1278_nl;
  mux_1280_nl <= MUX_s_1_2_2(or_3169_nl, or_3170_nl, fsm_output(1));
  GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c2 <= NOT(mux_1280_nl OR (fsm_output(8)));
  GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c3 <= and_dcpl_203 AND and_dcpl_237;
  and_601_nl <= (fsm_output(5)) AND (((CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")))
      AND (fsm_output(2))) OR (fsm_output(4)));
  mux_1283_nl <= MUX_s_1_2_2(and_1762_cse, and_601_nl, fsm_output(3));
  or_2203_nl <= nor_593_cse OR (fsm_output(4));
  mux_1282_nl <= MUX_s_1_2_2(mux_tmp_1281, or_2203_nl, fsm_output(0));
  nor_1060_nl <= NOT((fsm_output(3)) OR (fsm_output(5)) OR mux_1282_nl);
  mux_1284_nl <= MUX_s_1_2_2(mux_1283_nl, nor_1060_nl, fsm_output(6));
  GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c6 <= mux_1284_nl AND and_dcpl_295;
  attention_abs_qr_35_0_lpi_1_dfm_mx0c1 <= and_dcpl_192 AND and_dcpl_564 AND (NOT((fsm_output(7))
      OR (operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1(35))));
  nor_1102_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(1))) OR (fsm_output(8)) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR (NOT (fsm_output(6))));
  nor_1099_nl <= NOT((fsm_output(1)) OR (fsm_output(8)) OR (fsm_output(0)) OR (NOT
      (fsm_output(2))) OR (fsm_output(6)));
  nor_1100_nl <= NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(8))) OR (NOT LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4)
      OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(6)));
  mux_1401_nl <= MUX_s_1_2_2(nor_1099_nl, nor_1100_nl, fsm_output(3));
  nor_1101_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(1))) OR (fsm_output(8))
      OR (NOT (fsm_output(0))) OR (fsm_output(2)) OR (NOT (fsm_output(6))));
  mux_1402_nl <= MUX_s_1_2_2(mux_1401_nl, nor_1101_nl, fsm_output(7));
  and_1635_nl <= (fsm_output(5)) AND mux_1402_nl;
  RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c1 <= MUX_s_1_2_2(nor_1102_nl, and_1635_nl,
      fsm_output(4));
  mux_1407_nl <= MUX_s_1_2_2((NOT nor_tmp_285), and_1570_cse, fsm_output(5));
  mux_1408_nl <= MUX_s_1_2_2((NOT (fsm_output(5))), mux_1407_nl, fsm_output(3));
  mux_1409_nl <= MUX_s_1_2_2(mux_tmp_1027, mux_1408_nl, LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4);
  RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c4 <= (NOT mux_1409_nl) AND and_dcpl_413;
  mux_1447_nl <= MUX_s_1_2_2(or_270_cse, or_255_cse, and_1474_cse);
  and_1642_nl <= (fsm_output(6)) AND (fsm_output(3)) AND (NOT mux_1447_nl);
  mux_1444_nl <= MUX_s_1_2_2(and_dcpl_364, (fsm_output(4)), fsm_output(1));
  mux_1445_nl <= MUX_s_1_2_2((NOT mux_1444_nl), or_tmp_1221, fsm_output(0));
  mux_1442_nl <= MUX_s_1_2_2(or_tmp_11, mux_tmp_87, fsm_output(1));
  mux_1443_nl <= MUX_s_1_2_2(mux_1442_nl, mux_tmp_834, fsm_output(0));
  mux_1446_nl <= MUX_s_1_2_2(mux_1445_nl, mux_1443_nl, fsm_output(3));
  nor_1111_nl <= NOT((fsm_output(6)) OR mux_1446_nl);
  mux_1448_nl <= MUX_s_1_2_2(and_1642_nl, nor_1111_nl, fsm_output(7));
  CACHE_UPDATE_LOOP_3_k_2_0_sva_1_mx0c1 <= mux_1448_nl AND and_dcpl_1;
  nor_1118_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5)) OR (fsm_output(8)));
  nor_1119_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(0))) OR (fsm_output(6))
      OR (fsm_output(5)) OR (NOT (fsm_output(8))));
  mux_1464_nl <= MUX_s_1_2_2(nor_1118_nl, nor_1119_nl, fsm_output(4));
  and_1644_nl <= (NOT((fsm_output(1)) OR (NOT (fsm_output(3))))) AND mux_1464_nl;
  nor_1120_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(4)) OR (fsm_output(2))
      OR (fsm_output(0)) OR (fsm_output(6)) OR (NOT (fsm_output(5))) OR (fsm_output(8)));
  or_2363_nl <= (z_out_5(2)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(6))) OR
      (fsm_output(5)) OR (fsm_output(8));
  or_2362_nl <= (z_out_5(2)) OR (fsm_output(0)) OR (fsm_output(6)) OR (NOT (fsm_output(5)))
      OR (fsm_output(8));
  mux_1461_nl <= MUX_s_1_2_2(or_2363_nl, or_2362_nl, fsm_output(2));
  nor_1121_nl <= NOT((fsm_output(4)) OR mux_1461_nl);
  nor_1122_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(6))) OR (fsm_output(5))
      OR (fsm_output(8)));
  nor_1123_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(6)) OR (fsm_output(5))
      OR (fsm_output(8)));
  mux_1459_nl <= MUX_s_1_2_2(nor_1122_nl, nor_1123_nl, fsm_output(2));
  nor_1124_nl <= NOT((fsm_output(0)) OR CACHE_UPDATE_LOOP_1_and_tmp OR (fsm_output(6))
      OR (fsm_output(5)) OR (fsm_output(8)));
  nor_1125_nl <= NOT((z_out_5(2)) OR (NOT (fsm_output(0))) OR (fsm_output(6)) OR
      (fsm_output(5)) OR (fsm_output(8)));
  mux_1458_nl <= MUX_s_1_2_2(nor_1124_nl, nor_1125_nl, fsm_output(2));
  mux_1460_nl <= MUX_s_1_2_2(mux_1459_nl, mux_1458_nl, fsm_output(4));
  mux_1462_nl <= MUX_s_1_2_2(nor_1121_nl, mux_1460_nl, fsm_output(3));
  mux_1463_nl <= MUX_s_1_2_2(nor_1120_nl, mux_1462_nl, fsm_output(1));
  GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c1 <= MUX_s_1_2_2(and_1644_nl, mux_1463_nl,
      fsm_output(7));
  nor_1129_nl <= NOT((fsm_output(1)) OR RESHAPE_2D_TO_3D_LOOP_2_2_and_cse OR CONV_SL_1_1(fsm_output(8
      DOWNTO 4)/=STD_LOGIC_VECTOR'("01001")));
  nor_1130_nl <= NOT((NOT (fsm_output(1))) OR (NOT (z_out_5(2))) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 4)/=STD_LOGIC_VECTOR'("01100")));
  mux_1473_nl <= MUX_s_1_2_2(nor_1129_nl, nor_1130_nl, fsm_output(0));
  nor_1126_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 4)/=STD_LOGIC_VECTOR'("01001")));
  nor_1127_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT (fsm_output(4)))
      OR (fsm_output(8)));
  nor_1128_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(6)) OR (fsm_output(4))
      OR (fsm_output(8)));
  mux_1471_nl <= MUX_s_1_2_2(nor_1127_nl, nor_1128_nl, fsm_output(5));
  mux_1472_nl <= MUX_s_1_2_2(nor_1126_nl, mux_1471_nl, z_out_5(2));
  and_1646_nl <= nor_366_cse AND mux_1472_nl;
  mux_1474_nl <= MUX_s_1_2_2(mux_1473_nl, and_1646_nl, fsm_output(2));
  nor_1131_nl <= NOT((NOT (fsm_output(1))) OR (NOT CACHE_UPDATE_LOOP_1_and_tmp) OR
      CONV_SL_1_1(fsm_output(8 DOWNTO 4)/=STD_LOGIC_VECTOR'("01001")));
  nor_1132_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7)))
      OR (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1469_nl <= MUX_s_1_2_2(nor_1131_nl, nor_1132_nl, fsm_output(0));
  nor_1133_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR mux_1309_cse);
  nor_1134_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 4)/=STD_LOGIC_VECTOR'("01000")));
  mux_1467_nl <= MUX_s_1_2_2(nor_1133_nl, nor_1134_nl, fsm_output(1));
  nor_1135_nl <= NOT((NOT (fsm_output(1))) OR (NOT (z_out_5(2))) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 4)/=STD_LOGIC_VECTOR'("01001")));
  mux_1468_nl <= MUX_s_1_2_2(mux_1467_nl, nor_1135_nl, fsm_output(0));
  mux_1470_nl <= MUX_s_1_2_2(mux_1469_nl, mux_1468_nl, fsm_output(2));
  GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c2 <= MUX_s_1_2_2(mux_1474_nl, mux_1470_nl,
      fsm_output(3));
  or_2499_nl <= CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd) OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  mux_1586_nl <= MUX_s_1_2_2(nor_1026_cse, mux_tmp_1578, or_2499_nl);
  attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16_mx0c1 <= mux_1586_nl AND (NOT
      (fsm_output(8))) AND and_dcpl_814;
  nand_359_nl <= NOT(CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2=STD_LOGIC_VECTOR'("11"))
      AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd AND (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1));
  mux_1592_nl <= MUX_s_1_2_2(nor_1026_cse, mux_tmp_1578, nand_359_nl);
  attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16_mx0c1 <= mux_1592_nl AND (NOT
      (fsm_output(8))) AND and_dcpl_814;
  and_1811_cse <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  mux_2262_nl <= MUX_s_1_2_2(mux_tmp_1578, (NOT or_tmp_1354), and_1811_cse);
  mux_1594_nl <= MUX_s_1_2_2(mux_2262_nl, mux_tmp_1578, or_dcpl_332);
  attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16_mx0c1 <= mux_1594_nl AND (NOT
      (fsm_output(8))) AND and_dcpl_814;
  mux_1593_nl <= MUX_s_1_2_2(mux_tmp_1578, (NOT or_tmp_1354), and_1811_cse);
  mux_1595_nl <= MUX_s_1_2_2(mux_1593_nl, mux_tmp_1578, or_dcpl_342);
  attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16_mx0c1 <= mux_1595_nl AND (NOT
      (fsm_output(8))) AND and_dcpl_814;
  mux_1596_nl <= MUX_s_1_2_2(nor_1026_cse, mux_tmp_1578, or_2739_cse);
  attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16_mx0c1 <= mux_1596_nl AND (NOT
      (fsm_output(8))) AND and_dcpl_814;
  and_1659_nl <= (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(1)) AND
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  mux_1597_nl <= MUX_s_1_2_2(mux_tmp_1578, (NOT or_tmp_1354), and_1659_nl);
  mux_1598_nl <= MUX_s_1_2_2(mux_1597_nl, mux_tmp_1578, reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0));
  attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16_mx0c1 <= mux_1598_nl AND (NOT
      (fsm_output(8))) AND and_dcpl_814;
  mux_1599_nl <= MUX_s_1_2_2(nor_1026_cse, mux_tmp_1578, or_3039_cse);
  attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16_mx0c1 <= mux_1599_nl AND (NOT
      (fsm_output(8))) AND and_dcpl_814;
  nand_361_nl <= NOT(RESHAPE_2D_TO_3D_LOOP_2_2_and_cse AND (fsm_output(4)) AND (NOT
      (fsm_output(0))) AND (fsm_output(7)));
  nand_362_nl <= NOT((fsm_output(4)) AND (fsm_output(0)) AND (fsm_output(7)));
  mux_1605_nl <= MUX_s_1_2_2(nand_361_nl, nand_362_nl, fsm_output(3));
  nor_1160_nl <= NOT((fsm_output(2)) OR mux_1605_nl);
  nor_1161_nl <= NOT((NOT((fsm_output(3)) OR RESHAPE_2D_TO_3D_LOOP_2_2_and_cse))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (NOT (fsm_output(7))));
  nor_1162_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(0)) OR (NOT (fsm_output(7))));
  nor_1163_nl <= NOT((fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(7))));
  mux_1603_nl <= MUX_s_1_2_2(nor_1162_nl, nor_1163_nl, fsm_output(3));
  mux_1604_nl <= MUX_s_1_2_2(nor_1161_nl, mux_1603_nl, fsm_output(2));
  mux_1606_nl <= MUX_s_1_2_2(nor_1160_nl, mux_1604_nl, fsm_output(1));
  nor_1164_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(4))
      OR (fsm_output(0)) OR (NOT (fsm_output(7))));
  mux_1601_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), (fsm_output(7)), fsm_output(0));
  nor_1165_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("010"))
      OR mux_1601_nl);
  mux_1602_nl <= MUX_s_1_2_2(nor_1164_nl, nor_1165_nl, fsm_output(1));
  mux_1607_nl <= MUX_s_1_2_2(mux_1606_nl, mux_1602_nl, fsm_output(6));
  APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c0 <= mux_1607_nl AND and_dcpl_1;
  mux_1608_nl <= MUX_s_1_2_2(and_1555_cse, nor_749_cse, fsm_output(3));
  APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c2 <= mux_1608_nl AND and_dcpl_201
      AND and_dcpl_577 AND and_dcpl_45;
  and_1666_nl <= (fsm_output(4)) AND (NOT(nor_1106_cse OR (NOT (fsm_output(3))) OR
      (fsm_output(6))));
  nor_1169_nl <= NOT((CONV_SL_1_1(fsm_output(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111")))
      OR (fsm_output(6)));
  mux_1610_nl <= MUX_s_1_2_2(and_1666_nl, nor_1169_nl, fsm_output(5));
  and_1667_nl <= (fsm_output(8)) AND mux_1610_nl;
  nor_1170_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)));
  nor_1171_nl <= NOT((fsm_output(0)) OR (fsm_output(1)) OR (NOT (fsm_output(2)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))));
  mux_1609_nl <= MUX_s_1_2_2(nor_1170_nl, nor_1171_nl, fsm_output(4));
  and_1668_nl <= (NOT((fsm_output(8)) OR (NOT (fsm_output(5))))) AND mux_1609_nl;
  APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c3 <= MUX_s_1_2_2(and_1667_nl, and_1668_nl,
      fsm_output(7));
  or_2541_nl <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(4)));
  mux_1614_nl <= MUX_s_1_2_2(or_2541_nl, or_tmp_1392, fsm_output(6));
  or_3189_nl <= or_tmp_1392 OR (NOT (fsm_output(6)));
  mux_1615_nl <= MUX_s_1_2_2(mux_1614_nl, or_3189_nl, RESHAPE_2D_TO_3D_LOOP_2_2_and_cse);
  APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c4 <= (NOT mux_1615_nl) AND and_dcpl_226
      AND and_dcpl_885;
  apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c1 <= and_dcpl_732 AND
      and_dcpl_604;
  apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c8 <= and_dcpl_743 AND
      and_dcpl_551 AND and_dcpl_728;
  apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1 <= and_dcpl_732 AND
      and_dcpl_1000;
  attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c1 <= and_dcpl_732 AND and_dcpl_721;
  attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c6 <= and_dcpl_743 AND and_dcpl_552;
  attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0_mx0c1 <= and_dcpl_732 AND and_dcpl_591
      AND and_dcpl_462;
  or_2762_nl <= CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("11"))
      OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  mux_2060_nl <= MUX_s_1_2_2(nor_1026_cse, mux_tmp_1578, or_2762_nl);
  apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16_mx0c1 <= mux_2060_nl AND
      (NOT (fsm_output(8))) AND and_dcpl_814;
  or_2768_nl <= (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) OR CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd/=STD_LOGIC_VECTOR'("001"));
  mux_2069_nl <= MUX_s_1_2_2(or_1983_cse, mux_tmp_1562, or_2768_nl);
  apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16_mx0c1 <= (NOT(mux_2069_nl
      OR (fsm_output(8)))) AND and_dcpl_748;
  and_1781_cse <= (fsm_output(8)) AND (NOT(and_1782_cse OR CONV_SL_1_1(fsm_output(6
      DOWNTO 5)/=STD_LOGIC_VECTOR'("00"))));
  and_1778_nl <= ((CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      (z_out_5(2))) OR (fsm_output(5))) AND (fsm_output(6));
  mux_2138_nl <= MUX_s_1_2_2(and_1778_nl, (fsm_output(6)), fsm_output(2));
  or_1238_nl <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00"));
  mux_2136_nl <= MUX_s_1_2_2(or_1238_nl, (fsm_output(5)), or_3163_cse);
  mux_2137_nl <= MUX_s_1_2_2((fsm_output(6)), mux_2136_nl, nor_593_cse);
  mux_2139_cse <= MUX_s_1_2_2(mux_2138_nl, mux_2137_nl, fsm_output(3));
  or_2858_cse <= nor_305_cse OR (fsm_output(6));
  or_2856_cse <= nor_1026_cse OR (fsm_output(6));
  and_1780_nl <= (NOT(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 AND (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0))
      AND (fsm_output(0)) AND (fsm_output(5)))) AND (fsm_output(6));
  mux_2132_nl <= MUX_s_1_2_2(and_1780_nl, (fsm_output(6)), or_dcpl_672);
  mux_2133_nl <= MUX_s_1_2_2(or_2856_cse, mux_2132_nl, fsm_output(1));
  mux_2134_nl <= MUX_s_1_2_2(or_2858_cse, mux_2133_nl, fsm_output(2));
  mux_2135_nl <= MUX_s_1_2_2(mux_2134_nl, (fsm_output(6)), fsm_output(3));
  mux_2140_nl <= MUX_s_1_2_2(mux_2139_cse, mux_2135_nl, fsm_output(4));
  nor_1234_nl <= NOT((fsm_output(8)) OR (NOT mux_2140_nl));
  attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c1 <= MUX_s_1_2_2(and_1781_cse,
      nor_1234_nl, fsm_output(7));
  attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c9 <= and_dcpl_360 AND and_dcpl_355
      AND and_dcpl_539;
  attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx0c7 <= and_dcpl_360 AND and_dcpl_355
      AND and_dcpl_651;
  attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx0c7 <= and_dcpl_360 AND and_dcpl_355
      AND and_dcpl_656;
  and_1790_cse <= (NOT((fsm_output(0)) AND (fsm_output(5)))) AND (fsm_output(6));
  mux_2183_nl <= MUX_s_1_2_2(and_1790_cse, (fsm_output(6)), or_2671_cse);
  mux_2184_nl <= MUX_s_1_2_2(or_2856_cse, mux_2183_nl, fsm_output(1));
  mux_2185_nl <= MUX_s_1_2_2(or_2858_cse, mux_2184_nl, fsm_output(2));
  mux_2186_nl <= MUX_s_1_2_2(mux_2185_nl, (fsm_output(6)), fsm_output(3));
  mux_2191_nl <= MUX_s_1_2_2(mux_2139_cse, mux_2186_nl, fsm_output(4));
  nor_1261_nl <= NOT((fsm_output(8)) OR (NOT mux_2191_nl));
  attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c1 <= MUX_s_1_2_2(and_1781_cse,
      nor_1261_nl, fsm_output(7));
  attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c9 <= and_dcpl_360 AND and_dcpl_513
      AND and_dcpl_354;
  attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx0c7 <= and_dcpl_360 AND and_dcpl_513
      AND and_dcpl_458;
  attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx0c7 <= and_dcpl_360 AND and_dcpl_513
      AND and_dcpl_651;
  attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx0c7 <= and_dcpl_360 AND and_dcpl_513
      AND and_dcpl_656;
  mux_2211_nl <= MUX_s_1_2_2(and_1790_cse, (fsm_output(6)), or_2486_cse);
  mux_2212_nl <= MUX_s_1_2_2(or_2856_cse, mux_2211_nl, fsm_output(1));
  mux_2213_nl <= MUX_s_1_2_2(or_2858_cse, mux_2212_nl, fsm_output(2));
  mux_2214_nl <= MUX_s_1_2_2(mux_2213_nl, (fsm_output(6)), fsm_output(3));
  mux_2219_nl <= MUX_s_1_2_2(mux_2139_cse, mux_2214_nl, fsm_output(4));
  nor_1299_nl <= NOT((fsm_output(8)) OR (NOT mux_2219_nl));
  attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c1 <= MUX_s_1_2_2(and_1781_cse,
      nor_1299_nl, fsm_output(7));
  attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c9 <= and_dcpl_360 AND and_dcpl_355
      AND and_dcpl_512;
  attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx0c7 <= and_dcpl_360 AND and_dcpl_355
      AND and_dcpl_525;
  attention_abs_4_qr_35_0_lpi_1_dfm_mx0c1 <= and_dcpl_362 AND and_dcpl_198 AND CONV_SL_1_1(fsm_output(7
      DOWNTO 6)=STD_LOGIC_VECTOR'("11")) AND (NOT (operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1(35)));
  GEMM_3D_FLOAT_LOOP_4_l_and_ssc <= attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      AND (GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c0 OR GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c1
      OR GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c2 OR GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c3
      OR and_dcpl_193 OR and_dcpl_349 OR GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c6);
  GEMM_3D_FLOAT_LOOP_4_l_or_2_cse <= GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c1 OR
      and_dcpl_349;
  CACHE_UPDATE_LOOP_3_mux_3_nl <= MUX_v_40_16_2(attention_2_1_16_16_4_4_k_embed_0_0_0_sva_1,
      attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1, attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1,
      attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1, attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1,
      attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1, attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1,
      attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1,
      attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1,
      attention_2_1_16_16_4_4_k_embed_2_0_3_sva_1, attention_2_1_16_16_4_4_k_embed_3_0_0_sva_1,
      attention_2_1_16_16_4_4_k_embed_3_0_1_sva_1, attention_2_1_16_16_4_4_k_embed_3_0_2_sva_1,
      attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1, STD_LOGIC_VECTOR'( reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1));
  and_369_nl <= and_dcpl_322 AND and_dcpl_319 AND CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2=STD_LOGIC_VECTOR'("10"));
  attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d <= MUX_v_40_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_itm),40)),
      CACHE_UPDATE_LOOP_3_mux_3_nl, and_369_nl);
  TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_sdt_1(2
      DOWNTO 1)), 2), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1), 2), 3), 3));
  attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_nl),
      3)) & (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_sdt_1(0)) & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_pff <= and_dcpl_328;
  CACHE_UPDATE_LOOP_3_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(CACHE_UPDATE_LOOP_3_acc_sdt_1(2
      DOWNTO 1)), 2), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1), 2), 3), 3));
  attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(CACHE_UPDATE_LOOP_3_acc_nl),
      3)) & (CACHE_UPDATE_LOOP_3_acc_sdt_1(0)) & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_pff <= and_dcpl_318;
  CACHE_UPDATE_LOOP_3_1_mux_2_nl <= MUX_v_24_16_2(attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16, STD_LOGIC_VECTOR'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  CACHE_UPDATE_LOOP_3_1_CACHE_UPDATE_LOOP_3_1_mux_nl <= MUX_v_24_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_sdt(19
      DOWNTO 16)),24)), CACHE_UPDATE_LOOP_3_1_mux_2_nl, and_362_ssc);
  CACHE_UPDATE_LOOP_3_1_mux_3_nl <= MUX_v_16_16_2(attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0, STD_LOGIC_VECTOR'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  CACHE_UPDATE_LOOP_3_1_CACHE_UPDATE_LOOP_3_1_mux_1_nl <= MUX_v_16_2_2((CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_sdt(15
      DOWNTO 0)), CACHE_UPDATE_LOOP_3_1_mux_3_nl, and_362_ssc);
  attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d <= CACHE_UPDATE_LOOP_3_1_CACHE_UPDATE_LOOP_3_1_mux_nl
      & CACHE_UPDATE_LOOP_3_1_CACHE_UPDATE_LOOP_3_1_mux_1_nl;
  GEMM_3D_FLOAT_LOOP_4_1_acc_13_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(GEMM_3D_FLOAT_LOOP_4_1_acc_12_sdt_1(2
      DOWNTO 1)), 2), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1), 2), 3), 3));
  attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(GEMM_3D_FLOAT_LOOP_4_1_acc_13_nl),
      3)) & (GEMM_3D_FLOAT_LOOP_4_1_acc_12_sdt_1(0)) & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_pff <= and_dcpl_316;
  attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d <= GEMM_3D_FLOAT_LOOP_3_acc_6_tmp
      & (z_out_11(0)) & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1;
  GEMM_3D_FLOAT_LOOP_4_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(GEMM_3D_FLOAT_LOOP_4_acc_sdt_1(2
      DOWNTO 1)), 2), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1), 2), 3), 3));
  attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(GEMM_3D_FLOAT_LOOP_4_acc_nl),
      3)) & (GEMM_3D_FLOAT_LOOP_4_acc_sdt_1(0)) & (GEMM_3D_FLOAT_LOOP_4_acc_13_sdt_1(0))
      & (z_out_11(0));
  attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_pff <= and_dcpl_313;
  attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d <= TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_16_psp_1
      & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0)) & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_pff <= and_dcpl_289 AND and_dcpl_237;
  and_dcpl_1233 <= and_dcpl_222 AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd;
  and_dcpl_1248 <= CONV_SL_1_1(fsm_output(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"))
      AND and_dcpl_1 AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_1261 <= and_dcpl_61 AND (fsm_output(2)) AND (fsm_output(1)) AND (fsm_output(0))
      AND (fsm_output(3)) AND (NOT (fsm_output(5))) AND (NOT (fsm_output(6))) AND
      (fsm_output(7));
  nor_1345_nl <= NOT((fsm_output(6)) OR (fsm_output(2)) OR or_dcpl_959);
  nor_1346_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(2))) OR (fsm_output(4))
      OR (fsm_output(8)));
  mux_2299_nl <= MUX_s_1_2_2(nor_1345_nl, nor_1346_nl, fsm_output(7));
  and_dcpl_1273 <= mux_2299_nl AND (NOT (fsm_output(1))) AND (fsm_output(0)) AND
      (fsm_output(3)) AND (NOT (fsm_output(5)));
  and_dcpl_1294 <= nor_1314_cse AND (NOT (fsm_output(1))) AND (fsm_output(0)) AND
      (NOT (fsm_output(5))) AND (fsm_output(7));
  and_dcpl_1363 <= CONV_SL_1_1(fsm_output=STD_LOGIC_VECTOR'("011110101"));
  and_dcpl_1371 <= (NOT (fsm_output(8))) AND (fsm_output(4)) AND (NOT (fsm_output(1)))
      AND (fsm_output(2)) AND (NOT (fsm_output(0))) AND and_dcpl_198 AND CONV_SL_1_1(fsm_output(7
      DOWNTO 6)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_1379 <= and_dcpl_61 AND (fsm_output(1)) AND and_1555_cse AND and_dcpl_181
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_1385 <= (fsm_output(8)) AND (fsm_output(4)) AND (fsm_output(1)) AND and_1555_cse
      AND and_dcpl_181 AND nor_973_cse;
  and_dcpl_1391 <= and_dcpl_61 AND (fsm_output(1));
  and_dcpl_1392 <= and_dcpl_1391 AND nor_749_cse;
  and_dcpl_1393 <= and_dcpl_1392 AND and_dcpl_209;
  and_dcpl_1396 <= and_dcpl_201 AND (fsm_output(1));
  and_dcpl_1398 <= and_dcpl_1396 AND (NOT (fsm_output(2))) AND (fsm_output(0)) AND
      and_dcpl_209;
  and_dcpl_1401 <= (fsm_output(2)) AND (NOT (fsm_output(0)));
  and_dcpl_1403 <= and_dcpl_1396 AND and_dcpl_1401 AND (NOT (fsm_output(3))) AND
      (fsm_output(5)) AND nor_973_cse;
  and_dcpl_1406 <= and_dcpl_181 AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_1407 <= and_dcpl_1392 AND and_dcpl_1406;
  and_dcpl_1410 <= and_dcpl_1391 AND and_1555_cse AND and_dcpl_1406;
  and_dcpl_1415 <= and_dcpl_201 AND (NOT (fsm_output(1))) AND and_dcpl_1401 AND and_dcpl_198
      AND and_dcpl_45;
  nor_1378_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(2)));
  nor_1379_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(2))));
  mux_2288_nl <= MUX_s_1_2_2(nor_1378_nl, nor_1379_nl, fsm_output(6));
  and_dcpl_1420 <= mux_2288_nl AND and_dcpl_61 AND (fsm_output(1)) AND (fsm_output(0))
      AND (NOT (fsm_output(3))) AND (fsm_output(7));
  and_dcpl_1425 <= and_dcpl_61 AND (NOT (fsm_output(1))) AND and_1555_cse AND (fsm_output(3))
      AND (fsm_output(5)) AND and_dcpl_45;
  and_dcpl_1427 <= and_dcpl_181 AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_1429 <= and_dcpl_1391 AND and_dcpl_1401 AND and_dcpl_1427;
  and_dcpl_1431 <= and_dcpl_1396 AND and_1555_cse AND and_dcpl_1427;
  and_dcpl_1436 <= (fsm_output(8)) AND (fsm_output(4)) AND (fsm_output(1)) AND nor_749_cse
      AND and_dcpl_181 AND nor_973_cse;
  RMS_NORM_LOOP_1_1_or_3_ssc <= and_dcpl_1403 OR and_dcpl_1410 OR and_dcpl_1420 OR
      and_dcpl_1425 OR and_dcpl_1429;
  RMS_NORM_LOOP_1_1_or_1_ssc <= and_dcpl_1407 OR and_dcpl_1436;
  or_3261_nl <= (fsm_output(3)) OR nand_240_cse;
  or_3235_nl <= (fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(4));
  mux_2290_nl <= MUX_s_1_2_2(or_3235_nl, or_tmp_1128, fsm_output(0));
  mux_2291_nl <= MUX_s_1_2_2(mux_2290_nl, mux_1513_cse, fsm_output(3));
  mux_2292_nl <= MUX_s_1_2_2(or_3261_nl, mux_2291_nl, fsm_output(5));
  and_dcpl_1447 <= (NOT mux_2292_nl) AND and_dcpl_307 AND (fsm_output(7));
  RMS_NORM_LOOP_1_1_or_2_ssc <= and_dcpl_1407 OR and_dcpl_1425 OR and_dcpl_1429;
  and_1908_cse <= and_dcpl_61 AND (fsm_output(1)) AND (fsm_output(2)) AND (NOT (fsm_output(0)))
      AND (fsm_output(3)) AND (NOT (fsm_output(5))) AND (fsm_output(6)) AND (NOT
      (fsm_output(7)));
  mux_2266_nl <= MUX_s_1_2_2(nor_176_cse, and_1651_cse, fsm_output(2));
  nor_1348_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(1))) OR (fsm_output(4)));
  mux_2267_nl <= MUX_s_1_2_2(mux_2266_nl, nor_1348_nl, fsm_output(3));
  CACHE_UPDATE_LOOP_3_or_cse <= (mux_2267_nl AND (NOT (fsm_output(8))) AND (fsm_output(0))
      AND (NOT (fsm_output(5))) AND and_dcpl_45) OR and_1908_cse;
  nor_1350_nl <= NOT((fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(2)) OR (NOT
      and_1651_cse));
  mux_2268_nl <= MUX_s_1_2_2(nor_1053_cse, nor_1350_nl, fsm_output(7));
  nand_394_nl <= NOT((fsm_output(3)) AND (fsm_output(1)) AND (fsm_output(4)));
  mux_2270_nl <= MUX_s_1_2_2(nand_394_nl, or_tmp_704, fsm_output(5));
  CACHE_UPDATE_LOOP_3_or_1_cse <= (mux_2268_nl AND (NOT (fsm_output(8))) AND (fsm_output(3))
      AND (NOT (fsm_output(5)))) OR ((NOT(mux_2270_nl OR (fsm_output(8)))) AND (NOT
      (fsm_output(2))) AND (fsm_output(0)) AND and_dcpl_45);
  RMS_NORM_LOOP_1_1_or_5_cse <= and_dcpl_1398 OR and_dcpl_1403 OR and_dcpl_1431;
  RMS_NORM_LOOP_1_1_nor_seb <= NOT(and_dcpl_1398 OR and_dcpl_1431);
  RMS_NORM_LOOP_1_1_or_4_itm <= and_dcpl_1398 OR and_dcpl_1431;
  nand_398_nl <= NOT((fsm_output(1)) AND (fsm_output(4)));
  mux_2286_nl <= MUX_s_1_2_2(or_tmp_11, nand_398_nl, fsm_output(0));
  nor_1368_nl <= NOT((fsm_output(3)) OR mux_2286_nl);
  nor_1369_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011")));
  mux_2287_nl <= MUX_s_1_2_2(nor_1368_nl, nor_1369_nl, fsm_output(6));
  GEMM_3D_FLOAT_LOOP_1_or_ssc <= and_1908_cse OR (mux_2287_nl AND and_dcpl_1 AND
      (fsm_output(7)));
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        strm_out_rsci_idat_17_10 <= STD_LOGIC_VECTOR'( "00000000");
        strm_out_rsci_idat_9 <= '0';
        strm_out_rsci_idat_8 <= '0';
        strm_out_rsci_idat_7 <= '0';
        strm_out_rsci_idat_6 <= '0';
        strm_out_rsci_idat_5 <= '0';
        strm_out_rsci_idat_4 <= '0';
        strm_out_rsci_idat_3 <= '0';
        strm_out_rsci_idat_2 <= '0';
        strm_out_rsci_idat_31_18 <= STD_LOGIC_VECTOR'( "00000000000000");
      ELSIF ( for_1_for_and_cse = '1' ) THEN
        strm_out_rsci_idat_17_10 <= MUX_v_8_16_2((output_0_0_sva_2_15_0(15 DOWNTO
            8)), output_0_1_sva_2_15_8, (output_0_2_sva_2_15_0(15 DOWNTO 8)), (output_0_3_sva_2_15_0(15
            DOWNTO 8)), (output_0_4_sva_2_15_0(15 DOWNTO 8)), (output_0_5_sva_2_15_0(15
            DOWNTO 8)), (output_0_6_sva_2_15_0(15 DOWNTO 8)), (output_0_7_sva_2_15_0(15
            DOWNTO 8)), (output_0_8_sva_2_15_0(15 DOWNTO 8)), (output_0_9_sva_2_15_0(15
            DOWNTO 8)), (output_0_10_sva_2_15_0(15 DOWNTO 8)), (output_0_11_sva_2_15_0(15
            DOWNTO 8)), (output_0_12_sva_2_15_0(15 DOWNTO 8)), (output_0_13_sva_2_15_0(15
            DOWNTO 8)), (output_0_14_sva_2_15_0(15 DOWNTO 8)), (output_0_15_sva_2_15_0(15
            DOWNTO 8)), reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
        strm_out_rsci_idat_9 <= MUX_s_1_16_2((output_0_0_sva_2_15_0(7)), output_0_1_sva_2_7,
            (output_0_2_sva_2_15_0(7)), (output_0_3_sva_2_15_0(7)), (output_0_4_sva_2_15_0(7)),
            (output_0_5_sva_2_15_0(7)), (output_0_6_sva_2_15_0(7)), (output_0_7_sva_2_15_0(7)),
            (output_0_8_sva_2_15_0(7)), (output_0_9_sva_2_15_0(7)), (output_0_10_sva_2_15_0(7)),
            (output_0_11_sva_2_15_0(7)), (output_0_12_sva_2_15_0(7)), (output_0_13_sva_2_15_0(7)),
            (output_0_14_sva_2_15_0(7)), (output_0_15_sva_2_15_0(7)), reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
            & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
        strm_out_rsci_idat_8 <= MUX_s_1_16_2((output_0_0_sva_2_15_0(6)), output_0_1_sva_2_6,
            (output_0_2_sva_2_15_0(6)), (output_0_3_sva_2_15_0(6)), (output_0_4_sva_2_15_0(6)),
            (output_0_5_sva_2_15_0(6)), (output_0_6_sva_2_15_0(6)), (output_0_7_sva_2_15_0(6)),
            (output_0_8_sva_2_15_0(6)), (output_0_9_sva_2_15_0(6)), (output_0_10_sva_2_15_0(6)),
            (output_0_11_sva_2_15_0(6)), (output_0_12_sva_2_15_0(6)), (output_0_13_sva_2_15_0(6)),
            (output_0_14_sva_2_15_0(6)), (output_0_15_sva_2_15_0(6)), reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
            & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
        strm_out_rsci_idat_7 <= MUX_s_1_16_2((output_0_0_sva_2_15_0(5)), output_0_1_sva_2_5,
            (output_0_2_sva_2_15_0(5)), (output_0_3_sva_2_15_0(5)), (output_0_4_sva_2_15_0(5)),
            (output_0_5_sva_2_15_0(5)), (output_0_6_sva_2_15_0(5)), (output_0_7_sva_2_15_0(5)),
            (output_0_8_sva_2_15_0(5)), (output_0_9_sva_2_15_0(5)), (output_0_10_sva_2_15_0(5)),
            (output_0_11_sva_2_15_0(5)), (output_0_12_sva_2_15_0(5)), (output_0_13_sva_2_15_0(5)),
            (output_0_14_sva_2_15_0(5)), (output_0_15_sva_2_15_0(5)), reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
            & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
        strm_out_rsci_idat_6 <= MUX_s_1_16_2((output_0_0_sva_2_15_0(4)), output_0_1_sva_2_4,
            (output_0_2_sva_2_15_0(4)), (output_0_3_sva_2_15_0(4)), (output_0_4_sva_2_15_0(4)),
            (output_0_5_sva_2_15_0(4)), (output_0_6_sva_2_15_0(4)), (output_0_7_sva_2_15_0(4)),
            (output_0_8_sva_2_15_0(4)), (output_0_9_sva_2_15_0(4)), (output_0_10_sva_2_15_0(4)),
            (output_0_11_sva_2_15_0(4)), (output_0_12_sva_2_15_0(4)), (output_0_13_sva_2_15_0(4)),
            (output_0_14_sva_2_15_0(4)), (output_0_15_sva_2_15_0(4)), reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
            & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
        strm_out_rsci_idat_5 <= MUX_s_1_16_2((output_0_0_sva_2_15_0(3)), output_0_1_sva_2_3,
            (output_0_2_sva_2_15_0(3)), (output_0_3_sva_2_15_0(3)), (output_0_4_sva_2_15_0(3)),
            (output_0_5_sva_2_15_0(3)), (output_0_6_sva_2_15_0(3)), (output_0_7_sva_2_15_0(3)),
            (output_0_8_sva_2_15_0(3)), (output_0_9_sva_2_15_0(3)), (output_0_10_sva_2_15_0(3)),
            (output_0_11_sva_2_15_0(3)), (output_0_12_sva_2_15_0(3)), (output_0_13_sva_2_15_0(3)),
            (output_0_14_sva_2_15_0(3)), (output_0_15_sva_2_15_0(3)), reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
            & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
        strm_out_rsci_idat_4 <= MUX_s_1_16_2((output_0_0_sva_2_15_0(2)), output_0_1_sva_2_2,
            (output_0_2_sva_2_15_0(2)), (output_0_3_sva_2_15_0(2)), (output_0_4_sva_2_15_0(2)),
            (output_0_5_sva_2_15_0(2)), (output_0_6_sva_2_15_0(2)), (output_0_7_sva_2_15_0(2)),
            (output_0_8_sva_2_15_0(2)), (output_0_9_sva_2_15_0(2)), (output_0_10_sva_2_15_0(2)),
            (output_0_11_sva_2_15_0(2)), (output_0_12_sva_2_15_0(2)), (output_0_13_sva_2_15_0(2)),
            (output_0_14_sva_2_15_0(2)), (output_0_15_sva_2_15_0(2)), reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
            & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
        strm_out_rsci_idat_3 <= MUX_s_1_16_2((output_0_0_sva_2_15_0(1)), output_0_1_sva_2_1,
            (output_0_2_sva_2_15_0(1)), (output_0_3_sva_2_15_0(1)), (output_0_4_sva_2_15_0(1)),
            (output_0_5_sva_2_15_0(1)), (output_0_6_sva_2_15_0(1)), (output_0_7_sva_2_15_0(1)),
            (output_0_8_sva_2_15_0(1)), (output_0_9_sva_2_15_0(1)), (output_0_10_sva_2_15_0(1)),
            (output_0_11_sva_2_15_0(1)), (output_0_12_sva_2_15_0(1)), (output_0_13_sva_2_15_0(1)),
            (output_0_14_sva_2_15_0(1)), (output_0_15_sva_2_15_0(1)), reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
            & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
        strm_out_rsci_idat_2 <= MUX_s_1_16_2((output_0_0_sva_2_15_0(0)), output_0_1_sva_2_0,
            (output_0_2_sva_2_15_0(0)), (output_0_3_sva_2_15_0(0)), (output_0_4_sva_2_15_0(0)),
            (output_0_5_sva_2_15_0(0)), (output_0_6_sva_2_15_0(0)), (output_0_7_sva_2_15_0(0)),
            (output_0_8_sva_2_15_0(0)), (output_0_9_sva_2_15_0(0)), (output_0_10_sva_2_15_0(0)),
            (output_0_11_sva_2_15_0(0)), (output_0_12_sva_2_15_0(0)), (output_0_13_sva_2_15_0(0)),
            (output_0_14_sva_2_15_0(0)), (output_0_15_sva_2_15_0(0)), reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
            & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
        strm_out_rsci_idat_31_18 <= MUX_v_14_16_2(output_0_0_sva_2_29_16, output_0_1_sva_2_29_16,
            output_0_2_sva_2_29_16, output_0_3_sva_2_29_16, output_0_4_sva_2_29_16,
            output_0_5_sva_2_29_16, output_0_6_sva_2_29_16, output_0_7_sva_2_29_16,
            output_0_8_sva_2_29_16, output_0_9_sva_2_29_16, output_0_10_sva_2_29_16,
            output_0_11_sva_2_29_16, output_0_12_sva_2_29_16, output_0_13_sva_2_29_16,
            output_0_14_sva_2_29_16, output_0_15_sva_2_29_16, reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
            & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_39 <= '0';
        attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_38_0 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_3_0_0_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_attn_output_and_4_cse = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2 <= attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2_mx1;
        attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2 <= attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2_mx1;
        attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2 <= attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2_mx1;
        attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2 <= attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2_mx1;
        attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2 <= attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2_mx1;
        attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2 <= attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2_mx1;
        attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2 <= attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2_mx1;
        attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2 <= attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2_mx1;
        attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_39 <= attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_39;
        attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_38_0 <= attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_38_0;
        attention_2_1_16_16_4_4_attn_output_3_0_0_sva_2 <= MUX_v_40_2_2(acc_3_cse_40_1,
            attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3, nand_302_cse);
        attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2 <= attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2_mx1;
        attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2 <= attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2_mx1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_3_0_1_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (attention_2_1_16_16_4_4_attn_output_and_13_cse
          OR attention_2_1_16_16_4_4_attn_output_and_14_cse)) = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_3_0_1_sva_2 <= MUX_v_40_2_2(acc_3_cse_40_1,
            attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3, attention_2_1_16_16_4_4_attn_output_and_14_cse);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_3_0_2_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (attention_2_1_16_16_4_4_attn_output_and_15_cse
          OR attention_2_1_16_16_4_4_attn_output_and_16_cse)) = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_3_0_2_sva_2 <= MUX_v_40_2_2(acc_3_cse_40_1,
            attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3, attention_2_1_16_16_4_4_attn_output_and_16_cse);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_3_0_3_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (attention_2_1_16_16_4_4_attn_output_and_17_cse
          OR attention_2_1_16_16_4_4_attn_output_and_18_cse)) = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_3_0_3_sva_2 <= MUX_v_40_2_2(acc_3_cse_40_1,
            attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3, attention_2_1_16_16_4_4_attn_output_and_18_cse);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_attn_weights_and_36_cse = '1' ) THEN
        attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2_mx1,
            attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_3, and_dcpl_197);
        attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2_mx1,
            attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_3, and_dcpl_197);
        attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2_mx1,
            attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_3, and_dcpl_197);
        attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2_mx1,
            attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_3, and_dcpl_197);
        attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2_mx1,
            attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_3, and_dcpl_197);
        attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2_mx1,
            attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_3, and_dcpl_197);
        attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2_mx1,
            attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_3, and_dcpl_197);
        attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2_mx1,
            attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_3, and_dcpl_197);
        attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2_mx1,
            attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_3, and_dcpl_197);
        attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2_mx1,
            attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_3, and_dcpl_197);
        attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2_mx1,
            attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_3, and_dcpl_197);
        attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2_mx1,
            attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_3, and_dcpl_197);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_2_0_1_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_1_0_1_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_0_0_2_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_2_0_3_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_3_0_0_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_3_0_1_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_3_0_2_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_q_embed_and_5_cse = '1' ) THEN
        attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1 <= attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1_mx0w1;
        attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1 <= attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1_mx0w1;
        attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1 <= attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1_mx0w1;
        attention_2_1_16_16_4_4_q_embed_2_0_1_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
            attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1, or_dcpl_987);
        attention_2_1_16_16_4_4_q_embed_1_0_1_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
            attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1, or_dcpl_988);
        attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1 <= attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1_mx0w1;
        attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1 <= attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1_mx0w1;
        attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1 <= attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1_mx0w1;
        attention_2_1_16_16_4_4_q_embed_0_0_2_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
            attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1, or_dcpl_996);
        attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1 <= attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1_mx0w1;
        attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1 <= attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1_mx0w1;
        attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1 <= attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1_mx0w1;
        attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1 <= attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1_mx0w1;
        attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1 <= attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1_mx0w1;
        attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1 <= attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1_mx0w1;
        attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1 <= attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1_mx0w1;
        attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1 <= attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1_mx0w1;
        attention_2_1_16_16_4_4_k_embed_2_0_3_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
            attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3, or_dcpl_991);
        attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1 <= attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1_mx0w1;
        attention_2_1_16_16_4_4_k_embed_3_0_0_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
            attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3, or_dcpl_995);
        attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1 <= attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1_mx0w1;
        attention_2_1_16_16_4_4_k_embed_3_0_1_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
            attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3, or_dcpl_997);
        attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1 <= attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1_mx0w1;
        attention_2_1_16_16_4_4_k_embed_3_0_2_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
            attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3, or_dcpl_999);
        attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1 <= attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1_mx0w1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_embed_2_0_3_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_3_0_0_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_3_0_1_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_3_0_2_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_3_0_3_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd <= '0';
        reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd_1 <= '0';
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_47_40
            <= STD_LOGIC_VECTOR'( "00000000");
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_39
            <= '0';
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_38
            <= '0';
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_37
            <= '0';
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_36
            <= '0';
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_35
            <= '0';
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_34
            <= '0';
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_33
            <= '0';
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_32
            <= '0';
        operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_34 <= '0';
        operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_33_0 <= STD_LOGIC_VECTOR'(
            "0000000000000000000000000000000000");
        operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_39 <= '0';
        operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_38_35 <= STD_LOGIC_VECTOR'(
            "0000");
        SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_55 <= '0';
        SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_54_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000");
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_71_48
            <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_59_39
            <= STD_LOGIC_VECTOR'( "000000000000000000000");
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_38_0
            <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000");
        SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_39 <= '0';
        SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_38_0 <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000");
        reg_strm_out_rsci_iswt0_cse <= '0';
        reg_strm_in_rsci_iswt0_cse <= '0';
        reg_rms_norm_16_div_cmp_b_ftd_59_38 <= STD_LOGIC_VECTOR'( "0000000000000000000000");
        reg_rms_norm_16_div_cmp_b_ftd_37_0 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000");
        reg_rms_norm_16_div_cmp_b_ftd_1 <= '0';
        reg_rms_norm_16_div_cmp_a_ftd <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        reg_rms_norm_16_div_cmp_a_ftd_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        reg_rms_norm_16_div_cmp_a_ftd_1_7 <= '0';
        reg_rms_norm_16_div_cmp_a_ftd_1_6 <= '0';
        reg_rms_norm_16_div_cmp_a_ftd_1_5 <= '0';
        reg_rms_norm_16_div_cmp_a_ftd_1_4 <= '0';
        reg_rms_norm_16_div_cmp_a_ftd_1_3 <= '0';
        reg_rms_norm_16_div_cmp_a_ftd_1_2 <= '0';
        reg_rms_norm_16_div_cmp_a_ftd_1_1 <= '0';
        reg_rms_norm_16_div_cmp_a_ftd_1_0 <= '0';
        reg_RMS_NORM_LOOP_1_1_slc_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_mul_55_16_cse_1_slc
            <= STD_LOGIC_VECTOR'( "0000000000000000");
        operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_17_16
            <= STD_LOGIC_VECTOR'( "00");
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0 <= '0';
        attention_abs_3_qr_sva_38_0 <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000");
        RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_mux1h_itm <= '0';
        RMS_NORM_LOOP_2_and_29_ssc <= '0';
        RMS_NORM_LOOP_2_and_34_ssc <= '0';
        RMS_NORM_LOOP_2_and_30_m1c <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        reg_QUANTIZE_ACTIVATION_LOOP_3_quantized_value_slc_63_32_cse_slc <= STD_LOGIC_VECTOR'(
            "00000000");
        attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0 <= STD_LOGIC_VECTOR'(
            "0000000000000000");
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1 <= '0';
        LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000");
        APPLY_ROTARY_POS_EMB_LOOP_6_mul_3_itm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000");
        APPLY_ROTARY_POS_EMB_LOOP_6_mul_itm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000");
        APPLY_ROTARY_POS_EMB_LOOP_6_mul_1_itm <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000");
        TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_16_psp_1 <= STD_LOGIC_VECTOR'( "000");
        attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        operator_80_48_true_AC_TRN_AC_WRAP_operator_80_48_true_AC_TRN_AC_WRAP_slc_SOFTMAX_LOOP_4_sqr_56_1_itm_slc
            <= '0';
        attention_abs_5_qr_sva_38_0 <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000");
        attention_abs_7_qr_sva_38_0 <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000");
        RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_mux1h_itm <= '0';
        RMS_NORM_LOOP_2_2_and_29_ssc <= '0';
        RMS_NORM_LOOP_2_2_and_34_ssc <= '0';
        RMS_NORM_LOOP_2_2_and_30_m1c <= '0';
        output_0_7_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_7_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_8_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_8_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_6_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_6_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_9_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_9_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_5_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_5_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_10_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_10_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_4_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_4_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_11_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_11_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_3_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_3_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_12_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_12_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_2_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_2_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_13_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_13_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_1_lpi_3_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        output_0_1_lpi_3_7 <= '0';
        output_0_1_lpi_3_6 <= '0';
        output_0_1_lpi_3_5 <= '0';
        output_0_1_lpi_3_4 <= '0';
        output_0_1_lpi_3_3 <= '0';
        output_0_1_lpi_3_2 <= '0';
        output_0_1_lpi_3_1 <= '0';
        output_0_1_lpi_3_0 <= '0';
        output_0_14_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_14_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_0_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_0_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_15_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_15_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_15_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_0_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_14_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_1_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_13_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_2_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_12_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_3_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_11_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_4_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_10_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_5_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_9_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_6_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_8_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_7_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 = '1' ) THEN
        attention_2_1_16_16_4_4_q_embed_2_0_3_sva_1 <= attention_2_1_16_16_4_4_q_embed_mux_7_cse;
        attention_2_1_16_16_4_4_q_embed_3_0_0_sva_1 <= attention_2_1_16_16_4_4_q_embed_mux_9_cse;
        attention_2_1_16_16_4_4_q_embed_3_0_1_sva_1 <= attention_2_1_16_16_4_4_q_embed_mux_11_cse;
        attention_2_1_16_16_4_4_q_embed_3_0_2_sva_1 <= attention_2_1_16_16_4_4_q_embed_mux_13_cse;
        attention_2_1_16_16_4_4_q_embed_3_0_3_sva_1 <= attention_2_1_16_16_4_4_q_embed_mux_14_cse;
        reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd <= mux_816_ssc;
        reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd_1 <= NOT mux_816_ssc;
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_47_40
            <= MUX_v_8_2_2(STD_LOGIC_VECTOR'("00000000"), operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_nl,
            not_4947_nl);
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_39
            <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_1_nl AND (NOT or_dcpl_1048);
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_38
            <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_2_nl OR or_dcpl_1048;
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_37
            <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_3_nl OR or_dcpl_1048;
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_36
            <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_4_nl OR or_dcpl_1048;
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_35
            <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_5_nl OR or_dcpl_1048;
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_34
            <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_6_nl OR or_dcpl_1048;
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_33
            <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_7_nl OR or_dcpl_1048;
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_32
            <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_8_nl OR or_dcpl_1048;
        operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_34 <= MUX1HOT_s_1_7_2(compute_sqrt_guess_sva_34,
            attention_abs_qr_35_0_lpi_1_dfm_mx1_35, (compute_sqrt_for_acc_1_itm_40_1_1(34)),
            (attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_38_0(34)),
            (reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(34)), compute_sqrt_1_guess_sva_34,
            (compute_sqrt_1_for_acc_1_itm_40_1_1(34)), STD_LOGIC_VECTOR'( and_303_ssc
            & compute_sqrt_guess_or_1_ssc & and_dcpl_290 & and_dcpl_276 & and_dcpl_278
            & and_315_ssc & and_dcpl_292));
        operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_33_0 <= MUX1HOT_v_34_7_2(compute_sqrt_guess_sva_33_0,
            attention_abs_qr_35_0_lpi_1_dfm_mx1_34_1, (compute_sqrt_for_acc_1_itm_40_1_1(33
            DOWNTO 0)), (attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_38_0(33
            DOWNTO 0)), (reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(33 DOWNTO 0)), compute_sqrt_1_guess_sva_33_0,
            (compute_sqrt_1_for_acc_1_itm_40_1_1(33 DOWNTO 0)), STD_LOGIC_VECTOR'(
            and_303_ssc & compute_sqrt_guess_or_1_ssc & and_dcpl_290 & and_dcpl_276
            & and_dcpl_278 & and_315_ssc & and_dcpl_292));
        operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_39 <= rms_norm_16_mux1h_nl
            AND (NOT mux_851_ssc);
        operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_38_35 <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"),
            rms_norm_16_mux1h_9_nl, operator_40_24_true_AC_TRN_AC_WRAP_1_not_1_nl);
        SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_55 <= SOFTMAX_LOOP_5_mux_24_nl
            AND (NOT and_334_ssc);
        SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_54_16 <= MUX1HOT_v_39_3_2((SOFTMAX_LOOP_5_mux_12_psp_mx0w0(38
            DOWNTO 0)), reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1, STD_LOGIC_VECTOR'(
            "000000000000000000000010000000000000000"), STD_LOGIC_VECTOR'( and_dcpl_294
            & and_329_ssc & and_334_ssc));
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_71_48
            <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"), LINEAR_FORWARD_NO_MUL_LOOP_2_2_mux1h_2_nl,
            LINEAR_FORWARD_NO_MUL_LOOP_2_2_not_nl);
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_59_39
            <= MUX1HOT_v_21_5_2((z_out_9(59 DOWNTO 39)), (LINEAR_FORWARD_NO_MUL_LOOP_2_2_mul_mut(59
            DOWNTO 39)), STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_39,
            1),21)), STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd,
            1),21)), (LINEAR_FORWARD_NO_MUL_LOOP_2_3_mul_mut(59 DOWNTO 39)), STD_LOGIC_VECTOR'(
            LINEAR_FORWARD_NO_MUL_LOOP_2_2_or_1_cse & and_dcpl_260 & and_336_ssc
            & mux_856_ssc & and_dcpl_268));
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_38_0
            <= MUX1HOT_v_39_5_2((z_out_9(38 DOWNTO 0)), (LINEAR_FORWARD_NO_MUL_LOOP_2_2_mul_mut(38
            DOWNTO 0)), attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_38_0,
            reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1, (LINEAR_FORWARD_NO_MUL_LOOP_2_3_mul_mut(38
            DOWNTO 0)), STD_LOGIC_VECTOR'( LINEAR_FORWARD_NO_MUL_LOOP_2_2_or_1_cse
            & and_dcpl_260 & and_336_ssc & mux_856_ssc & and_dcpl_268));
        SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_39 <= MUX1HOT_s_1_3_2((softmax_1_4_3_sum_sva_1(39)),
            (compute_sqrt_1_for_acc_1_itm_40_1_1(39)), reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd,
            STD_LOGIC_VECTOR'( and_dcpl_304 & and_dcpl_292 & and_339_ssc));
        SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_38_0 <= MUX1HOT_v_39_3_2((softmax_1_4_3_sum_sva_1(38
            DOWNTO 0)), (compute_sqrt_1_for_acc_1_itm_40_1_1(38 DOWNTO 0)), reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1,
            STD_LOGIC_VECTOR'( and_dcpl_304 & and_dcpl_292 & and_339_ssc));
        reg_strm_out_rsci_iswt0_cse <= and_dcpl_306;
        reg_strm_in_rsci_iswt0_cse <= NOT(or_1851_cse OR (fsm_output(3)) OR or_1984_cse
            OR mux_862_nl OR or_255_cse);
        reg_rms_norm_16_div_cmp_b_ftd_59_38 <= MUX1HOT_v_22_5_2(STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(compute_sqrt_for_acc_1_itm_40_1_1(39),
            1),22)), STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd,
            1),22)), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2(60 DOWNTO 39)),
            (LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut(60 DOWNTO 39)), (LINEAR_FORWARD_NO_MUL_LOOP_2_mul_itm(59
            DOWNTO 38)), STD_LOGIC_VECTOR'( and_dcpl_290 & and_343_itm & and_dcpl_257
            & and_dcpl_260 & and_dcpl_310));
        reg_rms_norm_16_div_cmp_b_ftd_37_0 <= MUX1HOT_v_38_5_2((compute_sqrt_for_acc_1_itm_40_1_1(38
            DOWNTO 1)), (reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(38 DOWNTO 1)), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2(38
            DOWNTO 1)), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut(38 DOWNTO 1)), (LINEAR_FORWARD_NO_MUL_LOOP_2_mul_itm(37
            DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_290 & and_343_itm & and_dcpl_257
            & and_dcpl_260 & and_dcpl_310));
        reg_rms_norm_16_div_cmp_b_ftd_1 <= rms_norm_16_mux1h_10_nl AND (NOT and_dcpl_310);
        reg_rms_norm_16_div_cmp_a_ftd <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            rms_norm_16_mux1h_6_nl, rms_norm_16_not_nl);
        reg_rms_norm_16_div_cmp_a_ftd_1_15_8 <= MUX_v_8_2_2(STD_LOGIC_VECTOR'("00000000"),
            rms_norm_16_mux1h_7_nl, rms_norm_16_not_1_nl);
        reg_rms_norm_16_div_cmp_a_ftd_1_7 <= rms_norm_16_mux1h_11_nl AND (NOT rms_norm_16_div_cmp_a_mx0c0);
        reg_rms_norm_16_div_cmp_a_ftd_1_6 <= rms_norm_16_mux1h_13_nl AND (NOT rms_norm_16_div_cmp_a_mx0c0);
        reg_rms_norm_16_div_cmp_a_ftd_1_5 <= rms_norm_16_mux1h_14_nl AND (NOT rms_norm_16_div_cmp_a_mx0c0);
        reg_rms_norm_16_div_cmp_a_ftd_1_4 <= rms_norm_16_mux1h_15_nl AND (NOT rms_norm_16_div_cmp_a_mx0c0);
        reg_rms_norm_16_div_cmp_a_ftd_1_3 <= rms_norm_16_mux1h_16_nl AND (NOT rms_norm_16_div_cmp_a_mx0c0);
        reg_rms_norm_16_div_cmp_a_ftd_1_2 <= rms_norm_16_mux1h_17_nl AND (NOT rms_norm_16_div_cmp_a_mx0c0);
        reg_rms_norm_16_div_cmp_a_ftd_1_1 <= rms_norm_16_mux1h_18_nl AND (NOT rms_norm_16_div_cmp_a_mx0c0);
        reg_rms_norm_16_div_cmp_a_ftd_1_0 <= rms_norm_16_mux1h_19_nl OR rms_norm_16_div_cmp_a_mx0c0;
        reg_RMS_NORM_LOOP_1_1_slc_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_mul_55_16_cse_1_slc
            <= z_out_10(55 DOWNTO 40);
        operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_17_16
            <= operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z(17 DOWNTO 16);
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_15_8,
            attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8, and_dcpl_626);
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_7,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_38_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_6,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_39_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_5,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_40_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_4,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_41_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_3,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_42_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_2,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_43_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_1,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_44_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_0,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_15_8,
            attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8, and_dcpl_626);
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_1_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_7,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_24_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_6,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_5,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_26_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_4,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_27_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_3,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_28_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_2,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_29_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_1,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_30_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_0,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_15_8,
            attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8, and_dcpl_626);
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_2_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_7,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_10_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_6,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_11_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_5,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_12_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_4,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_13_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_3,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_14_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_2,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_15_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_1,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_16_nl,
            attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_0,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_15_8,
            attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8, and_dcpl_626);
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_3_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_7,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_17_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_6,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_18_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_5,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_19_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_4,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_20_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_3,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_21_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_2,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_22_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_1,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_23_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_0,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_15_8,
            attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8, and_dcpl_626);
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_4_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_7,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_31_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_6,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_32_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_5,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_33_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_4,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_34_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_3,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_35_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_2,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_36_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_1,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_37_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_0,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_15_8,
            attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8, and_dcpl_626);
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_5_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_7,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_45_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_6,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_46_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_5,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_47_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_4,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_48_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_3,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_49_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_2,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_50_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_1,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_51_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_0,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_15_8,
            attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8, and_dcpl_626);
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_6_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_7,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_52_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_6,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_53_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_5,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_54_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_4,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_55_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_3,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_56_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_2,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_57_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_1,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_58_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_0,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_15_8,
            attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8, and_dcpl_626);
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_7_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_7,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_59_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_6,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_60_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_5,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_61_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_4,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_62_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_3,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_63_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_2,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_64_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_1,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_65_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_0,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_15_8,
            attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8, and_dcpl_626);
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_8_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_7,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_66_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_6,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_67_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_5,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_68_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_4,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_69_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_3,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_70_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_2,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_71_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_1,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_72_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_0,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_15_8,
            attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8, and_dcpl_626);
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_9_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_7,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_73_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_6,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_74_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_5,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_75_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_4,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_76_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_3,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_77_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_2,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_78_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_1,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_79_nl,
            attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_0,
            STD_LOGIC_VECTOR'( and_dcpl_622 & and_dcpl_240 & and_dcpl_626));
        attention_abs_3_qr_sva_38_0 <= attention_abs_2_mux_2(38 DOWNTO 0);
        RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_mux1h_itm <= MUX1HOT_s_1_3_2((attention_abs_1_qr_sva_1(39)),
            reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1, (attention_abs_2_mux_2(39)),
            STD_LOGIC_VECTOR'( and_28_cse & RMS_NORM_LOOP_2_and_29_ssc_1 & RMS_NORM_LOOP_2_and_34_ssc_1));
        RMS_NORM_LOOP_2_and_29_ssc <= RMS_NORM_LOOP_2_and_29_ssc_1;
        RMS_NORM_LOOP_2_and_34_ssc <= RMS_NORM_LOOP_2_and_34_ssc_1;
        RMS_NORM_LOOP_2_and_30_m1c <= RMS_NORM_LOOP_2_and_30_m1c_1;
        attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_15_8,
            attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8, and_dcpl_626);
        reg_QUANTIZE_ACTIVATION_LOOP_3_quantized_value_slc_63_32_cse_slc <= z_out_10(63
            DOWNTO 56);
        attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_5_nl, not_4472_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_30_nl, not_4469_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_32_nl, not_4468_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_34_nl, not_4467_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_36_nl, not_4466_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_38_nl, not_4465_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_42_nl, not_4463_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_44_nl, not_4462_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_46_nl, not_4461_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_48_nl, not_4460_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_50_nl, not_4459_nl);
        apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            (attention_2_1_16_16_4_4_k_proj_re_mux1h_68_nl & attention_2_1_16_16_4_4_k_proj_re_mux1h_118_nl),
            not_4443_nl);
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_58_nl, not_4582_nl);
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_59_nl, not_4583_nl);
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_60_nl, not_4584_nl);
        attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_61_nl, not_4585_nl);
        attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_62_nl, not_4586_nl);
        attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_63_nl, not_4587_nl);
        attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_64_nl, not_4588_nl);
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_15_8,
            attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8, and_dcpl_626);
        LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1 <= (LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_2(1))
            AND (NOT mux_2100_ssc);
        LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0 <= QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_1_nl
            AND (NOT mux_2100_ssc);
        attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16 <= MUX_v_24_2_2(apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_39_16,
            attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16 <= MUX_v_24_2_2(LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48,
            attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16 <= MUX_v_24_2_2(apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_39_16,
            attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16 <= MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_39_16,
            attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16 <= MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16,
            attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_39_16,
            attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16 <= MUX_v_24_2_2(for_for_strm_in_tmp_sva_25_2,
            attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16,
            attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_39_16,
            attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_39_16,
            attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_39_16,
            attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16 <= MUX_v_24_2_2(apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16 <= MUX_v_24_2_2(apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_3_39_16,
            attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16 <= MUX_v_24_2_2(apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16 <= MUX_v_24_2_2(apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_3_39_16,
            attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16_mx1, and_dcpl_725);
        attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_39_16 <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16,
            attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16_mx0w1,
            attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16, STD_LOGIC_VECTOR'(
            and_dcpl_1073 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847));
        attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_39_16 <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16,
            attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16_mx0w1,
            attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16, STD_LOGIC_VECTOR'(
            and_dcpl_1073 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847));
        attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_39_16 <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16,
            attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16_mx0w1,
            attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16, STD_LOGIC_VECTOR'(
            and_dcpl_1073 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847));
        attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_39_16 <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16,
            attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16,
            attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16_mx0w1, STD_LOGIC_VECTOR'(
            operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse & and_dcpl_240 &
            attention_2_1_16_16_4_4_k_proj_re_or_17_cse & and_dcpl_207));
        attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_39_16 <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16,
            attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16_mx0w1,
            attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16, STD_LOGIC_VECTOR'(
            and_dcpl_1073 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847));
        APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm <= z_out_10(55 DOWNTO 0);
        APPLY_ROTARY_POS_EMB_LOOP_6_mul_3_itm <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'(
            CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(CONV_SIGNED(SIGNED((NOT and_dcpl_1363)
            & APPLY_ROTARY_POS_EMB_LOOP_6_mux_95_nl & APPLY_ROTARY_POS_EMB_LOOP_6_mux_96_nl
            & APPLY_ROTARY_POS_EMB_LOOP_6_APPLY_ROTARY_POS_EMB_LOOP_6_or_7_nl & APPLY_ROTARY_POS_EMB_LOOP_6_mux_97_nl
            & APPLY_ROTARY_POS_EMB_LOOP_6_mux_98_nl),16)), 16), 17) * SIGNED(APPLY_ROTARY_POS_EMB_LOOP_6_mux_99_nl
            & APPLY_ROTARY_POS_EMB_LOOP_6_mux_100_nl & APPLY_ROTARY_POS_EMB_LOOP_6_mux_101_nl)),
            56));
        APPLY_ROTARY_POS_EMB_LOOP_6_mul_itm <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'(
            SIGNED(LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48 & LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8
            & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1
            & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3
            & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5
            & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7)
            * SIGNED(reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd
            & reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1
            & reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2
            & (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3(7
            DOWNTO 5)) & '1' & (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3(4
            DOWNTO 0)))), 56));
        APPLY_ROTARY_POS_EMB_LOOP_6_mul_1_itm <= z_out_9(55 DOWNTO 0);
        TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_16_psp_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_15_sdt_1(2
            DOWNTO 1)), 2), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
            & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1), 2), 3), 3));
        attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2,
            attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_3,
            STD_LOGIC_VECTOR'( and_dcpl_1193 & and_dcpl_1194 & and_dcpl_1195));
        attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2,
            attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_3,
            STD_LOGIC_VECTOR'( and_dcpl_1193 & and_dcpl_1194 & and_dcpl_1195));
        attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2,
            attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_3,
            STD_LOGIC_VECTOR'( and_dcpl_1193 & and_dcpl_1194 & and_dcpl_1195));
        attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2,
            attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_3,
            STD_LOGIC_VECTOR'( and_dcpl_1193 & and_dcpl_1194 & and_dcpl_1195));
        attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2,
            attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_3,
            STD_LOGIC_VECTOR'( and_dcpl_1193 & and_dcpl_1194 & and_dcpl_1195));
        attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2,
            attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_3,
            STD_LOGIC_VECTOR'( and_dcpl_1193 & and_dcpl_1194 & and_dcpl_1195));
        attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2,
            attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_3,
            STD_LOGIC_VECTOR'( and_dcpl_1193 & and_dcpl_1194 & and_dcpl_1195));
        attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2,
            attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_3,
            STD_LOGIC_VECTOR'( and_dcpl_1193 & and_dcpl_1194 & and_dcpl_1195));
        attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2,
            attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_3,
            STD_LOGIC_VECTOR'( and_dcpl_1193 & and_dcpl_1194 & and_dcpl_1195));
        attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2,
            attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_3,
            STD_LOGIC_VECTOR'( and_dcpl_1193 & and_dcpl_1194 & and_dcpl_1195));
        attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2,
            attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_3,
            STD_LOGIC_VECTOR'( and_dcpl_1193 & and_dcpl_1194 & and_dcpl_1195));
        attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2,
            attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_3,
            STD_LOGIC_VECTOR'( and_dcpl_1193 & and_dcpl_1194 & and_dcpl_1195));
        operator_80_48_true_AC_TRN_AC_WRAP_operator_80_48_true_AC_TRN_AC_WRAP_slc_SOFTMAX_LOOP_4_sqr_56_1_itm_slc
            <= z_out_10(56);
        attention_abs_5_qr_sva_38_0 <= attention_abs_5_qr_sva_1(38 DOWNTO 0);
        attention_abs_7_qr_sva_38_0 <= attention_abs_6_mux_2(38 DOWNTO 0);
        RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_mux1h_itm <= MUX1HOT_s_1_3_2((attention_abs_5_qr_sva_1(39)),
            reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1, (attention_abs_6_mux_2(39)),
            STD_LOGIC_VECTOR'( RMS_NORM_LOOP_2_2_and_32_ssc_mx0w3 & RMS_NORM_LOOP_2_2_and_29_ssc_1
            & RMS_NORM_LOOP_2_2_and_34_ssc_1));
        RMS_NORM_LOOP_2_2_and_29_ssc <= RMS_NORM_LOOP_2_2_and_29_ssc_1;
        RMS_NORM_LOOP_2_2_and_34_ssc <= RMS_NORM_LOOP_2_2_and_34_ssc_1;
        RMS_NORM_LOOP_2_2_and_30_m1c <= RMS_NORM_LOOP_2_2_and_30_m1c_1;
        output_0_7_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_nl, not_4589_nl);
        output_0_7_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_44_nl, not_4590_nl);
        output_0_8_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_36_nl, not_4591_nl);
        output_0_8_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_45_nl, not_4592_nl);
        output_0_6_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_37_nl, not_4593_nl);
        output_0_6_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_46_nl, not_4594_nl);
        output_0_9_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_38_nl, not_4595_nl);
        output_0_9_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_47_nl, not_4596_nl);
        output_0_5_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_39_nl, not_4597_nl);
        output_0_5_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_48_nl, not_4598_nl);
        output_0_10_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_40_nl, not_4599_nl);
        output_0_10_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_49_nl, not_4600_nl);
        output_0_4_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_41_nl, not_4601_nl);
        output_0_4_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_50_nl, not_4602_nl);
        output_0_11_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_42_nl, not_4603_nl);
        output_0_11_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_51_nl, not_4604_nl);
        output_0_3_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_43_nl, not_4605_nl);
        output_0_3_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_52_nl, not_4606_nl);
        output_0_12_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_44_nl, not_4607_nl);
        output_0_12_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_53_nl, not_4608_nl);
        output_0_2_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_45_nl, not_4609_nl);
        output_0_2_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_54_nl, not_4610_nl);
        output_0_13_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_46_nl, not_4611_nl);
        output_0_13_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_55_nl, not_4612_nl);
        output_0_1_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_47_nl, not_4613_nl);
        output_0_1_lpi_3_15_8 <= MUX_v_8_2_2(STD_LOGIC_VECTOR'("00000000"), attention_2_1_16_16_4_4_k_proj_re_mux_56_nl,
            not_5055_nl);
        output_0_1_lpi_3_7 <= attention_2_1_16_16_4_4_k_proj_re_mux_60_nl AND (NOT
            and_dcpl_1154);
        output_0_1_lpi_3_6 <= attention_2_1_16_16_4_4_k_proj_re_mux_61_nl AND (NOT
            and_dcpl_1154);
        output_0_1_lpi_3_5 <= attention_2_1_16_16_4_4_k_proj_re_mux_62_nl AND (NOT
            and_dcpl_1154);
        output_0_1_lpi_3_4 <= attention_2_1_16_16_4_4_k_proj_re_mux_63_nl AND (NOT
            and_dcpl_1154);
        output_0_1_lpi_3_3 <= attention_2_1_16_16_4_4_k_proj_re_mux_64_nl AND (NOT
            and_dcpl_1154);
        output_0_1_lpi_3_2 <= attention_2_1_16_16_4_4_k_proj_re_mux_65_nl AND (NOT
            and_dcpl_1154);
        output_0_1_lpi_3_1 <= attention_2_1_16_16_4_4_k_proj_re_mux_66_nl AND (NOT
            and_dcpl_1154);
        output_0_1_lpi_3_0 <= attention_2_1_16_16_4_4_k_proj_re_mux_67_nl AND (NOT
            and_dcpl_1154);
        output_0_14_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_48_nl, not_4615_nl);
        output_0_14_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_57_nl, not_4616_nl);
        output_0_0_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_49_nl, not_4617_nl);
        output_0_0_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_58_nl, not_4618_nl);
        output_0_15_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_50_nl, not_4619_nl);
        output_0_15_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_59_nl, not_4620_nl);
        output_0_15_lpi_4_39_16 <= MUX_v_24_2_2(output_0_15_lpi_3_39_16, output_0_15_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_0_lpi_4_39_16 <= MUX_v_24_2_2(output_0_0_lpi_3_39_16, output_0_0_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_14_lpi_4_39_16 <= MUX_v_24_2_2(output_0_14_lpi_3_39_16, output_0_14_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_1_lpi_4_39_16 <= MUX_v_24_2_2(output_0_1_lpi_3_39_16, output_0_1_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_13_lpi_4_39_16 <= MUX_v_24_2_2(output_0_13_lpi_3_39_16, output_0_13_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_2_lpi_4_39_16 <= MUX_v_24_2_2(output_0_2_lpi_3_39_16, output_0_2_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_12_lpi_4_39_16 <= MUX_v_24_2_2(output_0_12_lpi_3_39_16, output_0_12_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_3_lpi_4_39_16 <= MUX_v_24_2_2(output_0_3_lpi_3_39_16, output_0_3_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_11_lpi_4_39_16 <= MUX_v_24_2_2(output_0_11_lpi_3_39_16, output_0_11_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_4_lpi_4_39_16 <= MUX_v_24_2_2(output_0_4_lpi_3_39_16, output_0_4_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_10_lpi_4_39_16 <= MUX_v_24_2_2(output_0_10_lpi_3_39_16, output_0_10_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_5_lpi_4_39_16 <= MUX_v_24_2_2(output_0_5_lpi_3_39_16, output_0_5_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_9_lpi_4_39_16 <= MUX_v_24_2_2(output_0_9_lpi_3_39_16, output_0_9_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_6_lpi_4_39_16 <= MUX_v_24_2_2(output_0_6_lpi_3_39_16, output_0_6_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_8_lpi_4_39_16 <= MUX_v_24_2_2(output_0_8_lpi_3_39_16, output_0_8_lpi_4_39_16_mx1,
            and_dcpl_1227);
        output_0_7_lpi_4_39_16 <= MUX_v_24_2_2(output_0_7_lpi_3_39_16, output_0_7_lpi_4_39_16_mx1,
            and_dcpl_1227);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_8 <= STD_LOGIC_VECTOR'(
            "00000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_7 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_6 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_5 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_4 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_3 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_2 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_1 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_0 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_13 <= STD_LOGIC_VECTOR'(
            "000");
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_12_8 <= STD_LOGIC_VECTOR'(
            "00000");
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_7 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_6 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_5 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_4 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_3 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_2 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_1 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_0 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_8 <= STD_LOGIC_VECTOR'(
            "00000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_7 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_6 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_5 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_4 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_3 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_2 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_1 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_0 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_8 <= STD_LOGIC_VECTOR'(
            "00000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_7 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_6 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_5 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_4 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_3 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_2 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_1 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_0 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_8 <= STD_LOGIC_VECTOR'(
            "00000000");
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd <=
            '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_1 <=
            '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_2 <=
            '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_3 <=
            '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_4 <=
            '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_5 <=
            '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_6 <=
            '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_7 <=
            '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_ftd <= STD_LOGIC_VECTOR'(
            "00000000");
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd <=
            '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_1 <=
            '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_2 <=
            '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_3 <=
            '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_4 <=
            '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_5 <=
            '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_6 <=
            '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_7 <=
            '0';
      ELSIF ( attention_2_1_16_16_4_4_v_proj_and_2_cse = '1' ) THEN
        attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_15_0 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
            attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0, or_dcpl_1010);
        attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_15_0 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
            attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0, or_dcpl_1012);
        attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_15_0 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
            attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0, or_dcpl_1014);
        attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_15_0 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
            attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0, or_dcpl_1016);
        attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_15_0 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
            attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0, or_dcpl_1018);
        attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0_mx0w1;
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16_mx0w1;
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_8 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_7 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_6 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_5 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_4 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_3 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_2 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_1 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_0 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16_mx0w1;
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_13 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_13;
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_12_8 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_12_8;
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_7 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_6 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_5 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_4 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_3 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_2 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_1 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_0 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16_mx0w1;
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_8 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_7 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_6 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_5 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_4 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_3 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_2 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_1 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_0 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_39_16 <= MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1,
            for_for_strm_in_tmp_sva_25_2, or_dcpl_1023);
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_8 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_7 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_6 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_5 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_4 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_3 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_2 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_1 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_0 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16 <= apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16_mx0w1;
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_8 <= apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd <=
            apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_1 <=
            apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_2 <=
            apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_3 <=
            apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_4 <=
            apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_5 <=
            apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_6 <=
            apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_7 <=
            apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16 <= apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16_mx0w1;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_ftd <= apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd <=
            apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_1 <=
            apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_2 <=
            apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_3 <=
            apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_4 <=
            apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_5 <=
            apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_6 <=
            apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
        reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_7 <=
            apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( apply_rotary_pos_emb_1_4_4_rotated_q_and_cse = '1' ) THEN
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2 <= MUX1HOT_v_40_7_2(apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm,
            apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2_mx0w1, attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1,
            attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2,
            GEMM_3D_FLOAT_LOOP_3_1_and_32_nl, attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2_mx1,
            STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_or_11_cse & and_dcpl_207
            & apply_rotary_pos_emb_1_4_4_rotated_q_or_12_cse & and_dcpl_204 & and_dcpl_220
            & and_dcpl_222 & and_dcpl_187));
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2 <= MUX1HOT_v_40_7_2(apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm,
            apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2_mx0w1, attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1,
            attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2,
            GEMM_3D_FLOAT_LOOP_3_1_and_34_nl, attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2_mx1,
            STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_or_11_cse & and_dcpl_207
            & apply_rotary_pos_emb_1_4_4_rotated_q_or_12_cse & and_dcpl_204 & and_dcpl_220
            & and_dcpl_222 & and_dcpl_187));
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2 <= MUX1HOT_v_40_7_2(apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm,
            apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2_mx0w1, attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1,
            attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2,
            GEMM_3D_FLOAT_LOOP_3_1_and_30_nl, attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2_mx1,
            STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_or_11_cse & and_dcpl_207
            & apply_rotary_pos_emb_1_4_4_rotated_q_or_12_cse & and_dcpl_204 & and_dcpl_220
            & and_dcpl_222 & and_dcpl_187));
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2 <= MUX1HOT_v_40_7_2(apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm,
            apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2_mx0w1, attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1,
            attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2,
            GEMM_3D_FLOAT_LOOP_3_1_and_40_nl, attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2_mx1,
            STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_or_11_cse & and_dcpl_207
            & apply_rotary_pos_emb_1_4_4_rotated_q_or_12_cse & and_dcpl_204 & and_dcpl_220
            & and_dcpl_222 & and_dcpl_187));
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2 <= MUX1HOT_v_40_7_2(apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm,
            apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2_mx0w1, attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1,
            attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2,
            GEMM_3D_FLOAT_LOOP_3_1_and_38_nl, attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2_mx1,
            STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_or_11_cse & and_dcpl_207
            & apply_rotary_pos_emb_1_4_4_rotated_q_or_12_cse & and_dcpl_204 & and_dcpl_220
            & and_dcpl_222 & and_dcpl_187));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT(mux_797_nl
          AND (NOT (fsm_output(8)))))) = '1' ) THEN
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2 <= MUX1HOT_v_40_6_2(apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w0,
            apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w3,
            attention_2_1_16_16_4_4_k_embed_0_0_0_sva_1, GEMM_3D_FLOAT_LOOP_3_1_and_42_nl,
            acc_3_cse_40_1, STD_LOGIC_VECTOR'( and_dcpl_207 & and_259_nl & and_dcpl_204
            & and_dcpl_216 & and_dcpl_222 & and_267_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1028)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_15 <= '0';
        attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_14_12 <= STD_LOGIC_VECTOR'( "000");
        attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_11_9 <= STD_LOGIC_VECTOR'( "000");
        attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_8 <= '0';
        attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_13 <= STD_LOGIC_VECTOR'( "000");
        attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0 <= STD_LOGIC_VECTOR'( "0000000000000");
        attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_ftd <= STD_LOGIC_VECTOR'(
            "00000000");
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd <= '0';
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_1 <= '0';
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_2 <= '0';
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_3 <= '0';
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_4 <= '0';
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_5 <= '0';
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_6 <= '0';
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_7 <= '0';
        attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd <= '0';
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_1 <= '0';
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_2 <= '0';
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_3 <= '0';
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_4 <= '0';
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_5 <= '0';
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_6 <= '0';
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_7 <= '0';
        attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_7 <= '0';
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_6 <= '0';
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_5 <= '0';
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_4 <= '0';
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_3 <= '0';
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_2 <= '0';
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_1 <= '0';
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_0 <= '0';
        attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_q_proj_and_23_cse = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_15_8;
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_7;
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_6;
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_5;
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_4;
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_3;
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_2;
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_1;
        attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_15_8;
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_7;
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_6;
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_5;
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_4;
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_3;
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_2;
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_1;
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_15_8;
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_7;
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_6;
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_5;
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_4;
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_3;
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_2;
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_1;
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_15_8;
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_7;
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_6;
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_5;
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_4;
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_3;
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_2;
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_1;
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_15_8;
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_7;
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_6;
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_5;
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_4;
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_3;
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_2;
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_1;
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_15_8;
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_7;
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_6;
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_5;
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_4;
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_3;
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_2;
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_1;
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_15_8;
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_7;
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_6;
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_5;
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_4;
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_3;
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_2;
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_1;
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_15_8;
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_7;
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_6;
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_5;
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_4;
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_3;
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_2;
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_1;
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_15 <= MUX_s_1_2_2((z_out(15)),
            operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_15,
            or_dcpl_1040);
        attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_14_12 <= MUX_v_3_2_2((z_out(14
            DOWNTO 12)), reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd,
            or_dcpl_1040);
        attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_11_9 <= MUX_v_3_2_2((z_out(11
            DOWNTO 9)), reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1,
            or_dcpl_1040);
        attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_8 <= MUX_s_1_2_2((z_out(8)), reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2,
            or_dcpl_1040);
        attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0 <= MUX_v_8_2_2((z_out(7 DOWNTO
            0)), reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3,
            or_dcpl_1040);
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_15_8;
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_7;
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_6;
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_5;
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_4;
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_3;
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_2;
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_1;
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0 <= attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_15_8;
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_7;
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_6;
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_5;
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_4;
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_3;
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_2;
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_1;
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0 <= attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_15_8;
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_7;
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_6;
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_5;
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_4;
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_3;
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_2;
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_1;
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_15_8;
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_7;
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_6;
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_5;
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_4;
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_3;
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_2;
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_1;
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_8 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_15_8;
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_7 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_7;
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_6 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_6;
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_5 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_5;
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_4 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_4;
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_3 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_3;
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_2 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_2;
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_1 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_1;
        attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_0 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_13 <= attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_15_13;
        attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0 <= attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0;
        attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_15_8 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_13_cse;
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_7 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_7;
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_6 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_6;
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_5 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_5;
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_4 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_4;
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_3 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_3;
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_2 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_2;
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_1 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_1;
        attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_0 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_0;
        attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16_mx0w1;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_ftd <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_15_8;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_7;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_1 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_6;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_2 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_5;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_3 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_4;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_4 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_3;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_5 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_2;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_6 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_1;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_7 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_8 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_15_8;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_7;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_1 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_6;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_2 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_5;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_3 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_4;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_4 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_3;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_5 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_2;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_6 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_1;
        reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_7 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_39_16 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
            for_for_strm_in_tmp_sva_25_2, or_dcpl_1017);
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_8 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_15_8;
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_7 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_7;
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_6 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_6;
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_5 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_5;
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_4 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_4;
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_3 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_3;
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_2 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_2;
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_1 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_1;
        attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_0 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_0;
        attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0_mx0w1;
        attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16_mx0w1;
        attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0_mx0w1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1030)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1031)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1033)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1035)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1037)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1038)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1039)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1040)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1041)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1042)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1043)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1044)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1045)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT or_dcpl_1046)
          AND and_dcpl_240) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        input_0_14_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_1_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_13_sva_1_39 <= '0';
        input_0_13_sva_1_38_0 <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000");
        input_0_2_sva_1_39 <= '0';
        input_0_2_sva_1_38_0 <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000");
        input_0_12_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_3_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_11_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_4_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_10_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_5_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_9_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_6_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_8_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_7_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( input_and_cse = '1' ) THEN
        input_0_14_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3,
            input_0_14_sva_2, and_dcpl_248);
        input_0_1_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3,
            input_0_1_sva_2, and_dcpl_248);
        input_0_13_sva_1_39 <= MUX_s_1_2_2(reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd,
            input_0_13_sva_2_39, and_dcpl_248);
        input_0_13_sva_1_38_0 <= MUX_v_39_2_2(reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1,
            input_0_13_sva_2_38_0, and_dcpl_248);
        input_0_2_sva_1_39 <= MUX_s_1_2_2(QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39,
            input_0_2_sva_2_39, and_dcpl_248);
        input_0_2_sva_1_38_0 <= MUX_v_39_2_2(QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0,
            input_0_2_sva_2_38_0, and_dcpl_248);
        input_0_12_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1,
            input_0_12_sva_2, and_dcpl_248);
        input_0_3_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3,
            input_0_3_sva_2, and_dcpl_248);
        input_0_11_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3,
            input_0_11_sva_2, and_dcpl_248);
        input_0_4_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3,
            input_0_4_sva_2, and_dcpl_248);
        input_0_10_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3,
            input_0_10_sva_2, and_dcpl_248);
        input_0_5_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3,
            input_0_5_sva_2, and_dcpl_248);
        input_0_9_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3,
            input_0_9_sva_2, and_dcpl_248);
        input_0_6_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3,
            input_0_6_sva_2, and_dcpl_248);
        input_0_8_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm, input_0_8_sva_2,
            and_dcpl_248);
        input_0_7_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1,
            input_0_7_sva_2, and_dcpl_248);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm <= STD_LOGIC_VECTOR'(
            "0000000000000000000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm <= STD_LOGIC_VECTOR'(
            "0000000000000000000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm <= STD_LOGIC_VECTOR'(
            "0000000000000000000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm <= STD_LOGIC_VECTOR'(
            "0000000000000000000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm <= STD_LOGIC_VECTOR'(
            "0000000000000000000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm <= STD_LOGIC_VECTOR'(
            "0000000000000000000000000000000000000000");
      ELSIF ( apply_rotary_pos_emb_1_4_4_rotated_q_and_3_cse = '1' ) THEN
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2_mx0w1;
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2_mx0w1;
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2_mx0w1;
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm <= apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2_mx0w1;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w0;
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm <= apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2_mx0w1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_15_8 <= STD_LOGIC_VECTOR'(
            "00000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_7 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_6 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_5 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_4 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_3 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_2 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_1 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_0 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd <= STD_LOGIC_VECTOR'(
            "00000000");
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_1 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_2 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_3 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_4 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_5 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_6 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_7 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_8 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( apply_rotary_pos_emb_1_4_4_rotated_k_and_6_cse = '1' ) THEN
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_15_8 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_7 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_6 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_5 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_4 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_2 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_1 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_0 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_1 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_2 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_4 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_5 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_6 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_7 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_8 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_39_16 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1;
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_39_16 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1;
        apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1;
        apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_15_8 <= STD_LOGIC_VECTOR'(
            "00000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_7 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_6 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_5 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_4 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_3 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_2 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_1 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_0 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd <= STD_LOGIC_VECTOR'(
            "00000000");
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_1 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_2 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_3 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_4 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_5 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_6 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_7 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_8 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( apply_rotary_pos_emb_1_4_4_rotated_k_and_7_cse = '1' ) THEN
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_15_8 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8;
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_7 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7;
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_6 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6;
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_5 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5;
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_4 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4;
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3;
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_2 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2;
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_1 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1;
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_0 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_1 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_2 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_4 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_5 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_6 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_7 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_8 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm;
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_39_16 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1;
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_39_16 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1;
        apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1;
        apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_15_8 <= STD_LOGIC_VECTOR'(
            "00000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_7 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_6 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_5 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_4 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_3 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_2 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_1 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_0 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd <= STD_LOGIC_VECTOR'(
            "00000000");
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_1 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_2 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_3 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_4 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_5 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_6 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_7 <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_8 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( apply_rotary_pos_emb_1_4_4_rotated_k_and_8_cse = '1' ) THEN
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_15_8 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8;
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_7 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7;
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_6 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6;
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_5 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5;
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_4 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4;
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3;
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_2 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2;
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_1 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1;
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_0 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_1 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_2 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_4 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_5 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_6 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_7 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm;
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_8 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm;
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_39_16 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1;
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_39_16 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1;
        apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1;
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (((NOT or_dcpl_1025)
          AND mux_902_nl) OR attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c0
          OR and_dcpl_344 OR and_dcpl_346 OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_349
          OR and_dcpl_351 OR attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c9))
          = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1 <= MUX1HOT_v_40_9_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),40)),
            input_0_0_sva_2, attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1, attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1_mx0w1,
            attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2, attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx2, (ATTN_2D_LOOP_3_mux_16_itm
            & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
            STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c0
            & and_dcpl_344 & and_dcpl_346 & and_dcpl_204 & and_dcpl_348 & and_dcpl_349
            & and_dcpl_351 & and_dcpl_352 & attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd <= '0';
        reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1 <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000");
      ELSIF ( GEMM_3D_FLOAT_LOOP_4_1_and_ssc = '1' ) THEN
        reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd <= rms_norm_16_variance_mux1h_nl AND
            GEMM_3D_FLOAT_LOOP_4_1_nand_itm;
        reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1 <= MUX_v_39_2_2(STD_LOGIC_VECTOR'("000000000000000000000000000000000000000"),
            rms_norm_16_variance_mux1h_1_nl, GEMM_3D_FLOAT_LOOP_4_1_nand_itm);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd <= '0';
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 <= '0';
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2 <= STD_LOGIC_VECTOR'(
            "00");
      ELSIF ( LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_ssc = '1' ) THEN
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd <= LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux_nl
            AND LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_5_itm;
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 <= LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_8_nl
            AND LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_5_itm;
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2 <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"),
            LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_9_nl, LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_5_itm);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd <= '0';
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 <= STD_LOGIC_VECTOR'(
            "00");
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 <= '0';
      ELSIF ( LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_and_ssc = '1' ) THEN
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd <= NOT((NOT(compute_sqrt_for_i_mux1h_nl
            AND (NOT LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c3))) OR LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c0);
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 <= NOT(MUX_v_2_2_2(compute_sqrt_for_i_nand_1_nl,
            STD_LOGIC_VECTOR'("11"), LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c0));
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 <= NOT((NOT(compute_sqrt_for_i_mux1h_2_nl
            OR LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c3)) OR LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        for_for_strm_in_tmp_sva_31_26 <= STD_LOGIC_VECTOR'( "000000");
        for_for_strm_in_tmp_sva_25_2 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( for_for_and_13_ssc = '1' ) THEN
        for_for_strm_in_tmp_sva_31_26 <= strm_in_rsci_idat_mxwt(29 DOWNTO 24);
        for_for_strm_in_tmp_sva_25_2 <= MUX_v_24_2_2((strm_in_rsci_idat_mxwt(23 DOWNTO
            0)), INIT_2D_MEM_LOOP_2_1_and_nl, for_for_strm_in_tmp_sva_31_2_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_1068)
          OR GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c0 OR GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c1
          OR GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c2 OR GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c4
          OR and_dcpl_313 OR GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c7 OR and_dcpl_316
          OR GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c9 OR GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c10)
          AND (mux_1063_nl OR (fsm_output(8)))) = '1' ) THEN
        GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm <= MUX1HOT_v_40_10_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),40)),
            input_0_8_sva_1, rms_norm_16_div_cmp_z_oreg, operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z,
            APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1, GEMM_3D_FLOAT_LOOP_4_mux_17_nl,
            STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SOFTMAX_LOOP_4_x_acc_2_nl), 40)),
            GEMM_3D_FLOAT_LOOP_4_1_mux_18_nl, z_out_2, (SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z(39
            DOWNTO 0)), STD_LOGIC_VECTOR'( GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c0
            & GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c1 & GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c2
            & GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c4 & and_dcpl_207 & and_dcpl_313
            & GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c7 & and_dcpl_316 & GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c9
            & GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39 <= '0';
        QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000000000000000000");
      ELSIF ( QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_and_ssc = '1' ) THEN
        QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39 <= MUX1HOT_s_1_13_2((strm_in_rsci_idat_mxwt(29)),
            input_0_2_sva_1_39, RMS_NORM_LOOP_2_mux_22_nl, QUANTIZE_ACTIVATION_LOOP_3_quantized_value_mux_nl,
            (APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1(39)), (attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d(39)),
            (attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1(39)), (attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1(39)),
            (attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1(39)), (attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1(39)),
            (SOFTMAX_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_cse_sva_1(39)),
            (attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d(39)), (z_out_2(39)), STD_LOGIC_VECTOR'(
            and_474_rgt & and_476_rgt & and_dcpl_438 & and_dcpl_439 & and_dcpl_374
            & and_480_rgt & for_for_and_14_rgt & for_for_and_15_rgt & for_for_and_16_rgt
            & for_for_and_17_rgt & and_485_rgt & and_486_rgt & for_for_or_1_rgt));
        QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0 <= MUX1HOT_v_39_13_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),39)),
            input_0_2_sva_1_38_0, RMS_NORM_LOOP_2_mux_24_nl, QUANTIZE_ACTIVATION_LOOP_3_quantized_value_mux_1_nl,
            (APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1(38 DOWNTO 0)), (attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d(38
            DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1(38 DOWNTO
            0)), (attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1(38 DOWNTO 0)),
            (attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1(38 DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1(38
            DOWNTO 0)), (SOFTMAX_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_cse_sva_1(38
            DOWNTO 0)), (attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d(38 DOWNTO 0)),
            (z_out_2(38 DOWNTO 0)), STD_LOGIC_VECTOR'( and_474_rgt & and_476_rgt
            & and_dcpl_438 & and_dcpl_439 & and_dcpl_374 & and_480_rgt & for_for_and_14_rgt
            & for_for_and_15_rgt & for_for_and_16_rgt & for_for_and_17_rgt & and_485_rgt
            & and_486_rgt & for_for_or_1_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_998)
          OR attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c0 OR attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c1
          OR (NOT mux_1079_itm) OR and_dcpl_204 OR and_dcpl_216 OR and_dcpl_348 OR
          and_dcpl_351 OR attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c7
          OR attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c9)) = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            for_for_mux1h_5_nl, attention_2_1_16_16_4_4_attn_output_2D_not_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_989)
          OR attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c0 OR attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c1
          OR and_dcpl_346 OR (NOT mux_1099_nl) OR and_dcpl_204 OR and_dcpl_348 OR
          and_dcpl_351 OR attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c7
          OR attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c9) AND (attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c0
          OR attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c1 OR and_dcpl_346
          OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_351 OR attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c7
          OR and_dcpl_352 OR attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c9))
          = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            for_for_mux1h_6_nl, attention_2_1_16_16_4_4_attn_output_2D_not_3_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd <= '0';
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000000000000000000");
      ELSIF ( apply_rotary_pos_emb_1_4_4_rotated_q_and_37_cse = '1' ) THEN
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd <= MUX1HOT_s_1_6_2((strm_in_rsci_idat_mxwt(29)),
            input_0_13_sva_1_39, (APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1(39)),
            attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_39, GEMM_3D_FLOAT_LOOP_3_1_and_36_nl,
            attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_39, STD_LOGIC_VECTOR'(
            apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c0 & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c1
            & and_dcpl_207 & and_dcpl_220 & and_dcpl_222 & and_dcpl_187));
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1 <= MUX1HOT_v_39_8_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),39)),
            input_0_13_sva_1_38_0, QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_dfm_1_38_0_1,
            QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_dfm_1_38_0_mx0w1, (APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1(38
            DOWNTO 0)), attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_38_0, GEMM_3D_FLOAT_LOOP_3_1_and_52_nl,
            attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_38_0, STD_LOGIC_VECTOR'(
            apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c0 & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c1
            & for_for_and_22_nl & and_dcpl_548 & and_dcpl_207 & and_dcpl_220 & and_dcpl_222
            & and_dcpl_187));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_attn_output_and_25_cse = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3 <= MUX1HOT_v_40_7_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),40)),
            input_0_1_sva_1, attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1, attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1_mx0w1,
            attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2, GEMM_3D_FLOAT_LOOP_3_1_and_28_nl,
            attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2_mx1, STD_LOGIC_VECTOR'(
            and_521_nl & and_523_nl & and_dcpl_346 & and_dcpl_204 & and_dcpl_220
            & and_dcpl_222 & and_dcpl_187));
        attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3 <= MUX1HOT_v_40_7_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),40)),
            input_0_14_sva_1, attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1, attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1_mx0w1,
            attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2, GEMM_3D_FLOAT_LOOP_3_1_and_29_nl,
            attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2_mx1, STD_LOGIC_VECTOR'(
            and_527_nl & and_529_nl & and_dcpl_346 & and_dcpl_204 & and_dcpl_220
            & and_dcpl_222 & and_dcpl_187));
        attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3 <= MUX1HOT_v_40_7_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),40)),
            input_0_6_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1_mx0w1,
            attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2, GEMM_3D_FLOAT_LOOP_3_1_and_31_nl,
            attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2_mx1, STD_LOGIC_VECTOR'(
            and_531_nl & and_533_nl & and_dcpl_346 & and_dcpl_204 & and_dcpl_220
            & and_dcpl_222 & and_dcpl_187));
        attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3 <= MUX1HOT_v_40_7_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),40)),
            input_0_9_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1_mx0w1,
            attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2, GEMM_3D_FLOAT_LOOP_3_1_and_33_nl,
            attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2_mx1, STD_LOGIC_VECTOR'(
            and_535_nl & and_537_nl & and_dcpl_346 & and_dcpl_204 & and_dcpl_220
            & and_dcpl_222 & and_dcpl_187));
        attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3 <= MUX1HOT_v_40_7_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),40)),
            input_0_5_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1_mx0w1,
            attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2, GEMM_3D_FLOAT_LOOP_3_1_and_35_nl,
            attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2_mx1, STD_LOGIC_VECTOR'(
            and_539_nl & and_541_nl & and_dcpl_346 & and_dcpl_204 & and_dcpl_220
            & and_dcpl_222 & and_dcpl_187));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_995)
          OR attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c0 OR attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c1
          OR and_dcpl_346 OR and_dcpl_204 OR attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c5
          OR and_dcpl_222 OR and_dcpl_187 OR attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c8
          OR attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c10) AND mux_1133_nl)
          = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            mux_nl, nor_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_997)
          OR attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c0 OR attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c1
          OR and_dcpl_346 OR (NOT mux_1147_itm) OR and_dcpl_204 OR and_dcpl_524 OR
          and_dcpl_222 OR and_dcpl_187 OR mux_tmp_1163 OR attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c10))
          = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            mux1h_nl, not_4622_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_999)
          OR attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c0 OR attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c1
          OR and_dcpl_346 OR (NOT mux_1177_itm) OR and_dcpl_204 OR and_dcpl_524 OR
          and_dcpl_222 OR and_dcpl_187 OR mux_tmp_1163 OR attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c10))
          = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            mux1h_1_nl, not_4624_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_1000)
          OR attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c0 OR attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c1
          OR and_dcpl_242 OR (NOT mux_1197_itm) OR and_dcpl_344 OR and_dcpl_346 OR
          and_dcpl_204 OR and_dcpl_524 OR and_dcpl_222 OR and_dcpl_187 OR attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c10
          OR attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c12)) = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            mux1h_2_nl, not_4626_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4 <= '0';
        LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_1_ssc = '1' ) THEN
        LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4 <= (LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_7_nl
            AND (NOT and_dcpl_477) AND LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_nand_seb)
            OR and_585_seb;
        LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0 <= MUX_v_4_2_2(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_4_nl,
            STD_LOGIC_VECTOR'("1111"), and_585_seb);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1 <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (and_dcpl_415
          OR and_dcpl_257)) = '1' ) THEN
        LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1 <= MUX_v_5_2_2(LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp,
            RMS_NORM_LOOP_2_2_acc_1_tmp, and_dcpl_257);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_abs_qr_35_0_lpi_1_dfm_35 <= '0';
        attention_abs_qr_35_0_lpi_1_dfm_34_0 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000");
      ELSIF ( attention_abs_qelse_and_ssc = '1' ) THEN
        attention_abs_qr_35_0_lpi_1_dfm_35 <= (attention_abs_qr_35_0_lpi_1_dfm_mx0w0(35))
            AND (NOT attention_abs_qr_35_0_lpi_1_dfm_mx0c1);
        attention_abs_qr_35_0_lpi_1_dfm_34_0 <= MUX_v_35_2_2((attention_abs_qr_35_0_lpi_1_dfm_mx0w0(34
            DOWNTO 0)), (operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1(34
            DOWNTO 0)), attention_abs_qr_35_0_lpi_1_dfm_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        compute_sqrt_guess_sva_34 <= '0';
        compute_sqrt_guess_sva_33_0 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000");
      ELSIF ( compute_sqrt_guess_and_ssc = '1' ) THEN
        compute_sqrt_guess_sva_34 <= MUX_s_1_2_2(attention_abs_qr_35_0_lpi_1_dfm_mx1_35,
            (compute_sqrt_for_acc_1_itm_40_1_1(34)), and_dcpl_290);
        compute_sqrt_guess_sva_33_0 <= MUX_v_34_2_2(attention_abs_qr_35_0_lpi_1_dfm_mx1_34_1,
            (compute_sqrt_for_acc_1_itm_40_1_1(33 DOWNTO 0)), and_dcpl_290);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_15
            <= '0';
        reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd
            <= STD_LOGIC_VECTOR'( "000");
        reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1
            <= STD_LOGIC_VECTOR'( "000");
        reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2
            <= '0';
      ELSIF ( operator_40_24_true_AC_TRN_AC_WRAP_1_and_ssc = '1' ) THEN
        operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_15
            <= MUX_s_1_2_2((operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z(15)),
            attention_2_1_16_16_4_4_q_proj_attention_2_1_16_16_4_4_q_proj_mux_12_nl,
            and_622_rgt);
        reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd
            <= MUX1HOT_v_3_4_2((operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z(14
            DOWNTO 12)), attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_14_12, (z_out(14
            DOWNTO 12)), (APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_itm(14
            DOWNTO 12)), STD_LOGIC_VECTOR'( and_615_itm & operator_40_24_true_AC_TRN_AC_WRAP_1_and_4_cse
            & and_1191_rgt & and_dcpl_583));
        reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1
            <= MUX1HOT_v_3_5_2((operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z(11
            DOWNTO 9)), (operator_40_24_true_AC_TRN_AC_WRAP_1_conc_1_itm_11_0(11
            DOWNTO 9)), attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_11_9, (z_out(11
            DOWNTO 9)), (APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_itm(11
            DOWNTO 9)), STD_LOGIC_VECTOR'( and_615_itm & and_dcpl_438 & operator_40_24_true_AC_TRN_AC_WRAP_1_and_4_cse
            & and_1191_rgt & and_dcpl_583));
        reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2
            <= MUX1HOT_s_1_6_2((operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z(8)),
            (operator_40_24_true_AC_TRN_AC_WRAP_1_conc_1_itm_11_0(8)), attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_8,
            (z_out(8)), (APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_itm(8)),
            (operator_40_24_true_AC_TRN_AC_WRAP_1_conc_3_itm_8_0(8)), STD_LOGIC_VECTOR'(
            and_615_itm & and_dcpl_438 & operator_40_24_true_AC_TRN_AC_WRAP_1_and_4_cse
            & and_1191_rgt & and_dcpl_583 & and_dcpl_448));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3
            <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( (operator_40_24_true_AC_TRN_AC_WRAP_1_and_ssc AND (NOT((NOT mux_1309_cse)
          AND and_dcpl_383 AND and_dcpl_338 AND and_dcpl_576))) = '1' ) THEN
        reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3
            <= MUX1HOT_v_8_8_2((operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z(7
            DOWNTO 0)), (operator_40_24_true_AC_TRN_AC_WRAP_1_conc_1_itm_11_0(7 DOWNTO
            0)), LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_itm,
            LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_itm,
            attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0, (z_out(7 DOWNTO 0)),
            (APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_itm(7
            DOWNTO 0)), (operator_40_24_true_AC_TRN_AC_WRAP_1_conc_3_itm_8_0(7 DOWNTO
            0)), STD_LOGIC_VECTOR'( and_615_itm & and_dcpl_438 & operator_40_24_true_AC_TRN_AC_WRAP_1_and_2_nl
            & and_dcpl_739 & operator_40_24_true_AC_TRN_AC_WRAP_1_and_4_cse & and_1191_rgt
            & and_dcpl_583 & and_dcpl_448));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_38_0 <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND and_dcpl_344)
          = '1' ) THEN
        QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_38_0 <= QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_dfm_1_38_0_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_quantized_hidden_states_0_9_sva_7 <= '0';
        reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_hidden_states_and_ssc = '1' ) THEN
        attention_2_1_16_16_4_4_quantized_hidden_states_0_9_sva_7 <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_cse;
        reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_quantized_hidden_states_0_6_sva_7 <= '0';
        reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_hidden_states_and_1_ssc = '1' ) THEN
        attention_2_1_16_16_4_4_quantized_hidden_states_0_6_sva_7 <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_cse;
        reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_quantized_hidden_states_0_8_sva_7 <= '0';
        reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_hidden_states_and_2_ssc = '1' ) THEN
        attention_2_1_16_16_4_4_quantized_hidden_states_0_8_sva_7 <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_cse;
        reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_quantized_hidden_states_0_7_sva_7 <= '0';
        reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_hidden_states_and_3_ssc = '1' ) THEN
        attention_2_1_16_16_4_4_quantized_hidden_states_0_7_sva_7 <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_cse;
        reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( RMS_NORM_LOOP_2_2_i_and_ssc = '1' ) THEN
        reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"),
            RMS_NORM_LOOP_2_2_i_mux1h_3_nl, RMS_NORM_LOOP_2_2_i_not_2_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 <= '0';
      ELSIF ( (RMS_NORM_LOOP_2_2_i_and_ssc AND (NOT(and_dcpl_1151 OR ((NOT and_dcpl_557)
          AND RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c4)))) = '1' ) THEN
        reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 <= RMS_NORM_LOOP_2_2_i_mux1h_6_nl
            AND (NOT RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        RMS_NORM_LOOP_2_2_i_4_0_sva_1 <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1434_nl
          OR (fsm_output(8)))) = '1' ) THEN
        RMS_NORM_LOOP_2_2_i_4_0_sva_1 <= MUX_v_5_2_2(RMS_NORM_LOOP_2_2_acc_1_tmp,
            LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp, and_dcpl_257);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1 <= '0';
        reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 <= '0';
      ELSIF ( CACHE_UPDATE_LOOP_3_k_and_ssc = '1' ) THEN
        reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1 <= MUX1HOT_s_1_3_2((z_out_3(2)), (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3(2)),
            (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(2)), STD_LOGIC_VECTOR'( and_dcpl_318
            & and_dcpl_328 & and_dcpl_635));
        reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 <= MUX1HOT_s_1_4_2(QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_3_nl,
            (z_out_3(1)), (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3(1)), (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(1)),
            STD_LOGIC_VECTOR'( CACHE_UPDATE_LOOP_3_k_2_0_sva_1_mx0c1 & and_dcpl_318
            & and_dcpl_328 & and_dcpl_635));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 <= '0';
      ELSIF ( (CACHE_UPDATE_LOOP_3_k_and_ssc AND (NOT(and_dcpl_629 OR compute_sqrt_for_i_and_2_cse)))
          = '1' ) THEN
        reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 <= MUX1HOT_s_1_6_2(RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_and_nl,
            QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_4_nl, (z_out_3(0)),
            (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3(0)), (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp(0)),
            (NOT QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1),
            STD_LOGIC_VECTOR'( CACHE_UPDATE_LOOP_3_k_and_1_nl & CACHE_UPDATE_LOOP_3_k_2_0_sva_1_mx0c1
            & and_dcpl_318 & and_dcpl_328 & and_dcpl_635 & and_dcpl_557));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd <= '0';
        reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 <= '0';
      ELSIF ( GEMM_3D_FLOAT_LOOP_1_i_and_ssc = '1' ) THEN
        reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd <= (z_out_5(1)) AND (NOT GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c2);
        reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 <= GEMM_3D_FLOAT_LOOP_1_i_mux_1_nl
            AND (NOT GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        input_0_0_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_1_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_2_sva_2_39 <= '0';
        input_0_2_sva_2_38_0 <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000");
        input_0_3_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_4_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_5_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_6_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_7_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_8_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_9_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_10_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_11_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_12_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_13_sva_2_39 <= '0';
        input_0_13_sva_2_38_0 <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000");
        input_0_14_sva_2 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        input_0_15_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( input_and_28_cse = '1' ) THEN
        input_0_0_sva_2 <= MUX_v_40_2_2((z_out_13_71_28(39 DOWNTO 0)), attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1,
            and_688_nl);
        input_0_1_sva_2 <= MUX_v_40_2_2((z_out_13_71_28(39 DOWNTO 0)), input_0_1_sva_1,
            and_693_nl);
        input_0_2_sva_2_39 <= MUX_s_1_2_2((z_out_13_71_28(39)), input_0_2_sva_1_39,
            and_699_ssc);
        input_0_2_sva_2_38_0 <= MUX_v_39_2_2((z_out_13_71_28(38 DOWNTO 0)), input_0_2_sva_1_38_0,
            and_699_ssc);
        input_0_3_sva_2 <= MUX_v_40_2_2((z_out_13_71_28(39 DOWNTO 0)), input_0_3_sva_1,
            and_704_nl);
        input_0_4_sva_2 <= MUX_v_40_2_2((z_out_13_71_28(39 DOWNTO 0)), input_0_4_sva_1,
            and_709_nl);
        input_0_5_sva_2 <= MUX_v_40_2_2((z_out_13_71_28(39 DOWNTO 0)), input_0_5_sva_1,
            and_713_nl);
        input_0_6_sva_2 <= MUX_v_40_2_2((z_out_13_71_28(39 DOWNTO 0)), input_0_6_sva_1,
            and_717_nl);
        input_0_7_sva_2 <= MUX_v_40_2_2((z_out_13_71_28(39 DOWNTO 0)), input_0_7_sva_1,
            and_721_nl);
        input_0_8_sva_2 <= MUX_v_40_2_2((z_out_13_71_28(39 DOWNTO 0)), input_0_8_sva_1,
            and_725_nl);
        input_0_9_sva_2 <= MUX_v_40_2_2((z_out_13_71_28(39 DOWNTO 0)), input_0_9_sva_1,
            and_729_nl);
        input_0_10_sva_2 <= MUX_v_40_2_2((z_out_13_71_28(39 DOWNTO 0)), input_0_10_sva_1,
            and_733_nl);
        input_0_11_sva_2 <= MUX_v_40_2_2((z_out_13_71_28(39 DOWNTO 0)), input_0_11_sva_1,
            and_737_nl);
        input_0_12_sva_2 <= MUX_v_40_2_2((z_out_13_71_28(39 DOWNTO 0)), input_0_12_sva_1,
            and_741_nl);
        input_0_13_sva_2_39 <= MUX_s_1_2_2((z_out_13_71_28(39)), input_0_13_sva_1_39,
            and_745_ssc);
        input_0_13_sva_2_38_0 <= MUX_v_39_2_2((z_out_13_71_28(38 DOWNTO 0)), input_0_13_sva_1_38_0,
            and_745_ssc);
        input_0_14_sva_2 <= MUX_v_40_2_2((z_out_13_71_28(39 DOWNTO 0)), input_0_14_sva_1,
            and_749_nl);
        input_0_15_sva_1 <= MUX_v_40_2_2((z_out_13_71_28(39 DOWNTO 0)), attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3,
            and_753_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva <= STD_LOGIC_VECTOR'(
            "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT(or_tmp_833
          OR nand_197_cse OR or_dcpl_1109 OR or_1984_cse))) = '1' ) THEN
        RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva <= z_out_13_71_28(39
            DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 <= '0';
      ELSIF ( APPLY_ROTARY_POS_EMB_LOOP_1_i_and_ssc = '1' ) THEN
        reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd <= (z_out_4(1)) AND mux_1512_itm;
        reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 <= APPLY_ROTARY_POS_EMB_LOOP_1_i_mux1h_5_nl
            AND mux_1512_itm;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd <= '0';
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_1 <= '0';
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_2 <= '0';
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_3 <= '0';
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_4 <= '0';
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_5 <= '0';
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_6 <= '0';
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_q_proj_and_4_ssc = '1' ) THEN
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1,
            attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_7,
            STD_LOGIC_VECTOR'( nor_1144_itm & and_dcpl_240 & and_dcpl_626));
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_1 <= MUX1HOT_s_1_3_2((NOT
            QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_6,
            attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_6, STD_LOGIC_VECTOR'( nor_1144_itm
            & and_dcpl_240 & and_dcpl_626));
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_2 <= MUX1HOT_s_1_3_2((NOT
            QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_5,
            attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_5, STD_LOGIC_VECTOR'( nor_1144_itm
            & and_dcpl_240 & and_dcpl_626));
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_3 <= MUX1HOT_s_1_3_2((NOT
            QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_4,
            attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_4, STD_LOGIC_VECTOR'( nor_1144_itm
            & and_dcpl_240 & and_dcpl_626));
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_4 <= MUX1HOT_s_1_3_2((NOT
            QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_3,
            attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_3, STD_LOGIC_VECTOR'( nor_1144_itm
            & and_dcpl_240 & and_dcpl_626));
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_5 <= MUX1HOT_s_1_3_2((NOT
            QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_2,
            attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_2, STD_LOGIC_VECTOR'( nor_1144_itm
            & and_dcpl_240 & and_dcpl_626));
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_6 <= MUX1HOT_s_1_3_2((NOT
            QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_1,
            attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_1, STD_LOGIC_VECTOR'( nor_1144_itm
            & and_dcpl_240 & and_dcpl_626));
        reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_7 <= MUX1HOT_s_1_3_2((NOT
            QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_0,
            attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_0, STD_LOGIC_VECTOR'( nor_1144_itm
            & and_dcpl_240 & and_dcpl_626));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_v_proj_re_and_cse = '1' ) THEN
        attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_4_nl, not_4557_nl);
        attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_8_nl, not_4558_nl);
        attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_12_nl, not_4559_nl);
        attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_16_nl, not_4560_nl);
        attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_20_nl, not_4561_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_21_nl, not_4562_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_q_proj_re_and_cse = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_35_nl, not_4441_nl);
        attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_34_nl, not_4440_nl);
        attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_33_nl, not_4439_nl);
        attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_32_nl, not_4438_nl);
        attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_31_nl, not_4437_nl);
        attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_30_nl, not_4436_nl);
        attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_29_nl, not_4435_nl);
        attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_28_nl, not_4434_nl);
        attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_27_nl, not_4433_nl);
        attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_26_nl, not_4432_nl);
        attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_25_nl, not_4431_nl);
        attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_24_nl, not_4430_nl);
        attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_23_nl, not_4429_nl);
        attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_22_nl, not_4428_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_7_sva_2_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_k_proj_re_and_1_cse = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_21_nl, not_4427_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_20_nl, not_4426_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_19_nl, not_4425_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_18_nl, not_4424_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_17_nl, not_4422_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux_16_nl, not_4415_nl);
        attention_2_1_16_16_4_4_k_proj_re_0_7_sva_2_39_16 <= MUX_v_24_2_2((rms_norm_16_div_cmp_z_oreg(39
            DOWNTO 16)), attention_2_1_16_16_4_4_k_proj_re_0_7_sva_1_39_16, and_1184_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (and_dcpl_619
          OR attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16_mx0c1 OR and_dcpl_843
          OR and_dcpl_207 OR and_dcpl_847)) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_40_nl, not_4423_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (and_dcpl_619
          OR attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16_mx0c1 OR and_dcpl_856
          OR and_dcpl_207 OR and_dcpl_847)) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_42_nl, not_4421_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (and_dcpl_619
          OR attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16_mx0c1 OR and_dcpl_860
          OR and_dcpl_207 OR and_dcpl_847)) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_43_nl, not_4420_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (and_dcpl_619
          OR attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16_mx0c1 OR and_dcpl_864
          OR and_dcpl_207 OR and_dcpl_847)) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_44_nl, not_4419_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (and_dcpl_619
          OR attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16_mx0c1 OR and_dcpl_868
          OR and_dcpl_207 OR and_dcpl_847)) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_45_nl, not_4418_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (and_dcpl_619
          OR attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16_mx0c1 OR and_dcpl_872
          OR and_dcpl_207 OR and_dcpl_847)) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_46_nl, not_4417_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (and_dcpl_619
          OR attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16_mx0c1 OR and_dcpl_876
          OR and_dcpl_207 OR and_dcpl_847)) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_47_nl, not_4416_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 <= '0';
      ELSIF ( APPLY_ROTARY_POS_EMB_LOOP_6_k_and_ssc = '1' ) THEN
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd <= GEMM_3D_FLOAT_LOOP_4_l_GEMM_3D_FLOAT_LOOP_4_l_mux_nl
            AND (NOT APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c0);
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 <= GEMM_3D_FLOAT_LOOP_4_l_mux1h_13_nl
            AND (NOT APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1641_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_26_nl, not_4471_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1644_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_28_nl, not_4470_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1727_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_40_nl, not_4464_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1816_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_43_nl, not_4458_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1825_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_42_nl, not_4457_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1834_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_41_nl, not_4456_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1843_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_40_nl, not_4455_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1852_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_39_nl, not_4454_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1861_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_38_nl, not_4453_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1870_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_37_nl, not_4452_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1878_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_36_nl, not_4451_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1887_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_35_nl, not_4450_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1896_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_34_nl, not_4449_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1905_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_33_nl, not_4448_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1914_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_32_nl, not_4447_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1923_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_31_nl, not_4446_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1932_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_30_nl, not_4445_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_1941_nl
          OR (fsm_output(8)))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux_29_nl, not_4444_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT((NOT mux_1946_nl)
          AND and_dcpl_259))) = '1' ) THEN
        attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_66_nl, not_4563_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT((NOT mux_1947_nl)
          AND and_dcpl_259))) = '1' ) THEN
        attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_67_nl, not_4564_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0 <= STD_LOGIC_VECTOR'(
            "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_1068)
          OR and_dcpl_619 OR apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c1
          OR and_dcpl_983 OR and_dcpl_240 OR and_dcpl_626 OR and_dcpl_739 OR apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c8)
          AND (NOT mux_1973_nl)) = '1' ) THEN
        apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            (attention_2_1_16_16_4_4_k_proj_re_mux1h_69_nl & attention_2_1_16_16_4_4_k_proj_re_mux1h_119_nl),
            not_4565_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_15_8 <= STD_LOGIC_VECTOR'(
            "00000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_7 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_6 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_5 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_4 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_3 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_2 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_1 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_0 <= '0';
      ELSIF ( apply_rotary_pos_emb_1_4_4_rotated_q_and_16_ssc = '1' ) THEN
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_15_8 <= MUX_v_8_2_2(STD_LOGIC_VECTOR'("00000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_70_nl, not_5074_nl);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_7 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_128_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_6 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_129_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_5 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_130_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_4 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_131_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_3 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_132_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_2 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_133_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_1 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_134_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_0 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_135_nl
            AND (NOT and_dcpl_619);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_8 <= STD_LOGIC_VECTOR'(
            "00000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_7 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_6 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_5 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_4 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_3 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_2 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_1 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_0 <= '0';
      ELSIF ( apply_rotary_pos_emb_1_4_4_rotated_q_and_17_ssc = '1' ) THEN
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_8 <= MUX_v_8_2_2(STD_LOGIC_VECTOR'("00000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_71_nl, not_5066_nl);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_7 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_120_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_6 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_121_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_5 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_122_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_4 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_123_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_3 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_124_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_2 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_125_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_1 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_126_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_0 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_127_nl
            AND (NOT and_dcpl_619);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_1145)
          OR and_dcpl_619 OR attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c1
          OR and_dcpl_410 OR and_dcpl_739 OR attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c6)
          AND mux_2012_nl) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_72_nl, not_4566_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT(or_dcpl_1146
          OR (NOT(mux_2022_nl OR (fsm_output(8)))))) OR and_dcpl_619 OR attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0_mx0c1
          OR and_dcpl_410)) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_73_nl, not_4567_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7 <= '0';
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6 <= '0';
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5 <= '0';
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4 <= '0';
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3 <= '0';
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2 <= '0';
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1 <= '0';
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0 <= '0';
      ELSIF ( APPLY_ROTARY_POS_EMB_LOOP_6_and_30_ssc = '1' ) THEN
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8 <= MUX_v_8_2_2(STD_LOGIC_VECTOR'("00000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_74_nl, not_5054_nl);
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_117_nl
            AND (NOT and_dcpl_619);
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_152_nl
            AND (NOT and_dcpl_619);
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_153_nl
            AND (NOT and_dcpl_619);
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_154_nl
            AND (NOT and_dcpl_619);
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_155_nl
            AND (NOT and_dcpl_619);
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_156_nl
            AND (NOT and_dcpl_619);
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_157_nl
            AND (NOT and_dcpl_619);
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_158_nl
            AND (NOT and_dcpl_619);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd <= STD_LOGIC_VECTOR'(
            "000");
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1 <= STD_LOGIC_VECTOR'(
            "0000000000000");
      ELSIF ( apply_rotary_pos_emb_1_4_4_rotated_q_and_18_ssc = '1' ) THEN
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_75_nl, not_4569_nl);
        reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1 <= MUX_v_13_2_2(STD_LOGIC_VECTOR'("0000000000000"),
            (attention_2_1_16_16_4_4_k_proj_re_mux1h_116_nl & attention_2_1_16_16_4_4_k_proj_re_mux1h_144_nl
            & attention_2_1_16_16_4_4_k_proj_re_mux1h_145_nl & attention_2_1_16_16_4_4_k_proj_re_mux1h_146_nl
            & attention_2_1_16_16_4_4_k_proj_re_mux1h_147_nl & attention_2_1_16_16_4_4_k_proj_re_mux1h_148_nl
            & attention_2_1_16_16_4_4_k_proj_re_mux1h_149_nl & attention_2_1_16_16_4_4_k_proj_re_mux1h_150_nl
            & attention_2_1_16_16_4_4_k_proj_re_mux1h_151_nl), not_5062_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_15_8 <= STD_LOGIC_VECTOR'(
            "00000000");
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_7 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_6 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_5 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_4 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_3 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_2 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_1 <= '0';
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_0 <= '0';
      ELSIF ( apply_rotary_pos_emb_1_4_4_rotated_q_and_19_ssc = '1' ) THEN
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_15_8 <= MUX_v_8_2_2(STD_LOGIC_VECTOR'("00000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_76_nl, not_5088_nl);
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_7 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_136_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_6 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_137_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_5 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_138_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_4 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_139_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_3 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_140_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_2 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_141_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_1 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_142_nl
            AND (NOT and_dcpl_619);
        apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_0 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_143_nl
            AND (NOT and_dcpl_619);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT((NOT mux_2038_nl)
          AND and_dcpl_259))) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_77_nl, not_4571_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT((NOT mux_2039_nl)
          AND and_dcpl_259))) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_78_nl, not_4572_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT((NOT mux_2040_nl)
          AND and_dcpl_259))) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_79_nl, not_4573_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_2051_nl
          OR (fsm_output(7)))) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_80_nl, not_4574_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT((NOT mux_2052_nl)
          AND and_dcpl_259))) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_81_nl, not_4575_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT((NOT mux_2053_nl)
          AND and_dcpl_259))) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_82_nl, not_4576_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT((NOT mux_2054_nl)
          AND and_dcpl_259))) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_83_nl, not_4577_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT((NOT mux_2055_nl)
          AND and_dcpl_259))) = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_15_0 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            attention_2_1_16_16_4_4_k_proj_re_mux1h_84_nl, not_4578_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (mux_2059_nl
          OR (fsm_output(8)))) = '1' ) THEN
        apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_51_nl, not_4414_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT(or_dcpl_1068
          OR (NOT(mux_2063_nl OR (fsm_output(8)))))) OR and_dcpl_619 OR apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16_mx0c1
          OR and_dcpl_1003)) = '1' ) THEN
        apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_52_nl, not_4413_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT((NOT mux_2068_nl)
          AND and_dcpl_581))) = '1' ) THEN
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_53_nl, not_4412_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT(or_dcpl_1068
          OR ((NOT mux_tmp_2067) AND and_dcpl_581))) OR and_dcpl_619 OR apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16_mx0c1
          OR and_dcpl_959)) = '1' ) THEN
        apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_54_nl, not_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT(or_dcpl_1145
          OR and_dcpl_1055)) OR and_dcpl_619 OR and_dcpl_726 OR and_dcpl_410)) =
          '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_55_nl, not_4579_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (and_dcpl_619
          OR and_dcpl_726 OR and_dcpl_257 OR and_dcpl_1033 OR and_dcpl_983 OR and_dcpl_240
          OR and_dcpl_1034 OR and_dcpl_207 OR and_dcpl_213 OR and_dcpl_583 OR and_dcpl_265))
          = '1' ) THEN
        LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_56_nl, not_4580_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (and_dcpl_619
          OR and_dcpl_726 OR and_dcpl_257 OR and_dcpl_1011 OR and_dcpl_983 OR and_dcpl_240
          OR and_dcpl_207 OR and_dcpl_847 OR and_dcpl_583)) = '1' ) THEN
        APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16 <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
            attention_2_1_16_16_4_4_v_proj_re_mux1h_57_nl, not_4581_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_7 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_6 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_5 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_4 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_3 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_2 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_1 <= '0';
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_0 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_q_proj_and_5_ssc = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_7 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_nl,
            attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_7,
            STD_LOGIC_VECTOR'( nor_1228_ssc & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_6 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse,
            attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_6,
            STD_LOGIC_VECTOR'( nor_1228_ssc & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_5 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse,
            attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_5,
            STD_LOGIC_VECTOR'( nor_1228_ssc & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_4 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse,
            attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_4,
            STD_LOGIC_VECTOR'( nor_1228_ssc & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_3 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse,
            attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_3,
            STD_LOGIC_VECTOR'( nor_1228_ssc & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_2 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse,
            attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_2,
            STD_LOGIC_VECTOR'( nor_1228_ssc & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_1 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse,
            attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_1,
            STD_LOGIC_VECTOR'( nor_1228_ssc & and_dcpl_240 & and_dcpl_626));
        attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_0 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse,
            attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_0,
            STD_LOGIC_VECTOR'( nor_1228_ssc & and_dcpl_240 & and_dcpl_626));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd <= STD_LOGIC_VECTOR'(
            "00000000");
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd <= STD_LOGIC_VECTOR'(
            "00000000");
      ELSIF ( APPLY_ROTARY_POS_EMB_LOOP_6_and_28_cse = '1' ) THEN
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd <= MUX1HOT_v_8_6_2((drf_output_sdt_2_sva_15_0_mx0w0(15
            DOWNTO 8)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_8, attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_15_8,
            apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8,
            apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_8, APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_nl,
            STD_LOGIC_VECTOR'( and_dcpl_257 & and_dcpl_1073 & and_dcpl_240 & and_dcpl_207
            & and_dcpl_847 & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd <= MUX1HOT_v_8_6_2((z_out(15
            DOWNTO 8)), attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_8, attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_15_8,
            apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8,
            apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_8, APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_nl,
            STD_LOGIC_VECTOR'( and_dcpl_257 & and_dcpl_1073 & and_dcpl_240 & and_dcpl_207
            & and_dcpl_847 & and_dcpl_583));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1 <= '0';
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0 <= '0';
      ELSIF ( APPLY_ROTARY_POS_EMB_LOOP_6_and_31_cse = '1' ) THEN
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm(7)),
            (drf_output_sdt_2_sva_15_0_mx0w0(7)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_7,
            attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_7, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7,
            apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_7, APPLY_ROTARY_POS_EMB_LOOP_6_mux_66_nl,
            STD_LOGIC_VECTOR'( and_dcpl_888 & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240
            & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm(6)),
            (drf_output_sdt_2_sva_15_0_mx0w0(6)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_6,
            attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_6, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6,
            apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_6, APPLY_ROTARY_POS_EMB_LOOP_6_mux_74_nl,
            STD_LOGIC_VECTOR'( and_dcpl_888 & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240
            & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm(5)),
            (drf_output_sdt_2_sva_15_0_mx0w0(5)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_5,
            attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_5, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5,
            apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_5, APPLY_ROTARY_POS_EMB_LOOP_6_mux_75_nl,
            STD_LOGIC_VECTOR'( and_dcpl_888 & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240
            & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm(4)),
            (drf_output_sdt_2_sva_15_0_mx0w0(4)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_4,
            attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_4, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4,
            apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_4, APPLY_ROTARY_POS_EMB_LOOP_6_mux_76_nl,
            STD_LOGIC_VECTOR'( and_dcpl_888 & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240
            & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm(3)),
            (drf_output_sdt_2_sva_15_0_mx0w0(3)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_3,
            attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_3, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3,
            apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_3, APPLY_ROTARY_POS_EMB_LOOP_6_mux_77_nl,
            STD_LOGIC_VECTOR'( and_dcpl_888 & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240
            & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm(2)),
            (drf_output_sdt_2_sva_15_0_mx0w0(2)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_2,
            attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_2, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2,
            apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_2, APPLY_ROTARY_POS_EMB_LOOP_6_mux_78_nl,
            STD_LOGIC_VECTOR'( and_dcpl_888 & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240
            & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm(1)),
            (drf_output_sdt_2_sva_15_0_mx0w0(1)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_1,
            attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_1, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1,
            apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_1, APPLY_ROTARY_POS_EMB_LOOP_6_mux_79_nl,
            STD_LOGIC_VECTOR'( and_dcpl_888 & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240
            & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm(0)),
            (drf_output_sdt_2_sva_15_0_mx0w0(0)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_0,
            attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_0, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0,
            apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_0, APPLY_ROTARY_POS_EMB_LOOP_6_mux_80_nl,
            STD_LOGIC_VECTOR'( and_dcpl_888 & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240
            & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm(7)),
            (z_out(7)), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd,
            attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_7, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7,
            reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_61_nl, STD_LOGIC_VECTOR'( and_dcpl_888
            & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847
            & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm(6)),
            (z_out(6)), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_1,
            attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_6, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6,
            reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_1,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_81_nl, STD_LOGIC_VECTOR'( and_dcpl_888
            & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847
            & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm(5)),
            (z_out(5)), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_2,
            attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_5, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5,
            reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_2,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_82_nl, STD_LOGIC_VECTOR'( and_dcpl_888
            & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847
            & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm(4)),
            (z_out(4)), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_3,
            attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_4, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4,
            reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_3,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_83_nl, STD_LOGIC_VECTOR'( and_dcpl_888
            & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847
            & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm(3)),
            (z_out(3)), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_4,
            attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_3, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3,
            reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_4,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_84_nl, STD_LOGIC_VECTOR'( and_dcpl_888
            & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847
            & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm(2)),
            (z_out(2)), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_5,
            attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_2, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2,
            reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_5,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_85_nl, STD_LOGIC_VECTOR'( and_dcpl_888
            & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847
            & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm(1)),
            (z_out(1)), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_6,
            attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_1, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1,
            reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_6,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_86_nl, STD_LOGIC_VECTOR'( and_dcpl_888
            & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847
            & and_dcpl_583));
        reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm(0)),
            (z_out(0)), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_7,
            attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_0, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0,
            reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_7,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_87_nl, STD_LOGIC_VECTOR'( and_dcpl_888
            & and_dcpl_257 & and_dcpl_1073 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847
            & and_dcpl_583));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_re_0_0_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_14_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_13_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_12_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_11_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_4_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_10_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_5_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_9_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_6_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_8_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_7_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_q_proj_re_0_15_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_q_proj_re_and_29_cse = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_re_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_14_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_13_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_12_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_11_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_4_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_10_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_5_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_9_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_6_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_8_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_7_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_q_proj_re_0_15_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16_mx1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_proj_re_0_15_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_0_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_14_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_13_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_12_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_11_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_4_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_10_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_5_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_9_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_6_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_8_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_k_proj_re_0_7_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_k_proj_re_and_65_cse = '1' ) THEN
        attention_2_1_16_16_4_4_k_proj_re_0_15_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_14_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_13_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_12_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_11_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_4_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_10_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_5_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_9_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_6_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_8_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_k_proj_re_0_7_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16_mx1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_v_proj_re_0_15_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_0_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_14_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_13_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_12_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_4_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_10_sva_1_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_5_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_9_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_6_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_8_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_7_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_v_proj_re_and_32_cse = '1' ) THEN
        attention_2_1_16_16_4_4_v_proj_re_0_15_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_14_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_13_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_12_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_4_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_10_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_5_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_9_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_6_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_8_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16_mx1;
        attention_2_1_16_16_4_4_v_proj_re_0_7_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16_mx1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        LINEAR_FORWARD_NO_MUL_LOOP_2_mul_itm <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000000000000000000000000");
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_mul_mut <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000000000000000000000000");
        LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000");
      ELSIF ( LINEAR_FORWARD_NO_MUL_LOOP_2_and_cse = '1' ) THEN
        LINEAR_FORWARD_NO_MUL_LOOP_2_mul_itm <= z_out_10(59 DOWNTO 0);
        LINEAR_FORWARD_NO_MUL_LOOP_2_2_mul_mut <= z_out_9;
        LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut <= LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd <= '0';
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1 <= '0';
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2 <= '0';
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3 <= '0';
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4 <= '0';
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5 <= '0';
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6 <= '0';
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7 <= '0';
      ELSIF ( LINEAR_FORWARD_NO_MUL_LOOP_2_1_and_29_ssc = '1' ) THEN
        LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8 <= MUX1HOT_v_8_7_2((z_out_1(15
            DOWNTO 8)), attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_15_8, RESHAPE_2D_TO_3D_LOOP_3_1_mux_13_cse,
            apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_8, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8,
            (APPLY_ROTARY_POS_EMB_LOOP_6_mux_32_nl & APPLY_ROTARY_POS_EMB_LOOP_6_mux_70_nl
            & APPLY_ROTARY_POS_EMB_LOOP_6_mux_71_nl & APPLY_ROTARY_POS_EMB_LOOP_6_mux_72_nl),
            (drf_output_sdt_3_sva_15_0_mx0w3(15 DOWNTO 8)), STD_LOGIC_VECTOR'( and_dcpl_257
            & operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse & and_dcpl_240
            & attention_2_1_16_16_4_4_k_proj_re_or_17_cse & and_dcpl_207 & and_dcpl_583
            & and_dcpl_265));
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd <= MUX1HOT_s_1_7_2((z_out_1(7)),
            attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_7, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_7,
            apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_7, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_50_nl, (drf_output_sdt_3_sva_15_0_mx0w3(7)),
            STD_LOGIC_VECTOR'( and_dcpl_257 & operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse
            & and_dcpl_240 & attention_2_1_16_16_4_4_k_proj_re_or_17_cse & and_dcpl_207
            & and_dcpl_583 & and_dcpl_265));
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1 <= MUX1HOT_s_1_7_2((z_out_1(6)),
            attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_6, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_6,
            apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_6, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_51_nl, (drf_output_sdt_3_sva_15_0_mx0w3(6)),
            STD_LOGIC_VECTOR'( and_dcpl_257 & operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse
            & and_dcpl_240 & attention_2_1_16_16_4_4_k_proj_re_or_17_cse & and_dcpl_207
            & and_dcpl_583 & and_dcpl_265));
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2 <= MUX1HOT_s_1_7_2((z_out_1(5)),
            attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_5, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_5,
            apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_5, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_52_nl, (drf_output_sdt_3_sva_15_0_mx0w3(5)),
            STD_LOGIC_VECTOR'( and_dcpl_257 & operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse
            & and_dcpl_240 & attention_2_1_16_16_4_4_k_proj_re_or_17_cse & and_dcpl_207
            & and_dcpl_583 & and_dcpl_265));
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3 <= MUX1HOT_s_1_7_2((z_out_1(4)),
            attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_4, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_4,
            apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_4, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_53_nl, (drf_output_sdt_3_sva_15_0_mx0w3(4)),
            STD_LOGIC_VECTOR'( and_dcpl_257 & operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse
            & and_dcpl_240 & attention_2_1_16_16_4_4_k_proj_re_or_17_cse & and_dcpl_207
            & and_dcpl_583 & and_dcpl_265));
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4 <= MUX1HOT_s_1_7_2((z_out_1(3)),
            attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_3, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_3,
            apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_3, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_54_nl, (drf_output_sdt_3_sva_15_0_mx0w3(3)),
            STD_LOGIC_VECTOR'( and_dcpl_257 & operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse
            & and_dcpl_240 & attention_2_1_16_16_4_4_k_proj_re_or_17_cse & and_dcpl_207
            & and_dcpl_583 & and_dcpl_265));
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5 <= MUX1HOT_s_1_7_2((z_out_1(2)),
            attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_2, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_2,
            apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_2, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_55_nl, (drf_output_sdt_3_sva_15_0_mx0w3(2)),
            STD_LOGIC_VECTOR'( and_dcpl_257 & operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse
            & and_dcpl_240 & attention_2_1_16_16_4_4_k_proj_re_or_17_cse & and_dcpl_207
            & and_dcpl_583 & and_dcpl_265));
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6 <= MUX1HOT_s_1_7_2((z_out_1(1)),
            attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_1, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_1,
            apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_1, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_56_nl, (drf_output_sdt_3_sva_15_0_mx0w3(1)),
            STD_LOGIC_VECTOR'( and_dcpl_257 & operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse
            & and_dcpl_240 & attention_2_1_16_16_4_4_k_proj_re_or_17_cse & and_dcpl_207
            & and_dcpl_583 & and_dcpl_265));
        reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7 <= MUX1HOT_s_1_7_2((z_out_1(0)),
            attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_0, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_0,
            apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_0, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0,
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_57_nl, (drf_output_sdt_3_sva_15_0_mx0w3(0)),
            STD_LOGIC_VECTOR'( and_dcpl_257 & operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse
            & and_dcpl_240 & attention_2_1_16_16_4_4_k_proj_re_or_17_cse & and_dcpl_207
            & and_dcpl_583 & and_dcpl_265));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_39_16 <= STD_LOGIC_VECTOR'(
            "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_7 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_6 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_5 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_4 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_3 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_2 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_1 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_0 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_15_13 <= STD_LOGIC_VECTOR'(
            "000");
        attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0 <= STD_LOGIC_VECTOR'( "0000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_7 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_6 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_5 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_4 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_3 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_2 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_1 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_0 <= '0';
        attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_v_proj_re_and_95_cse = '1' ) THEN
        attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_0_sva_1_39_16, and_dcpl_1084);
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_1_sva_1_39_16, and_dcpl_1088);
        attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_2_sva_1_39_16, and_dcpl_1091);
        attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_3_sva_1_39_16, and_dcpl_1094);
        attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_4_sva_1_39_16, and_dcpl_1097);
        attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_5_sva_1_39_16, and_dcpl_1100);
        attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_6_sva_1_39_16, and_dcpl_1103);
        attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_7_sva_1_39_16, and_dcpl_1106);
        attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_8_sva_1_39_16, and_dcpl_1109);
        attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_9_sva_1_39_16, and_dcpl_1112);
        attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_10_sva_1_39_16, and_dcpl_1115);
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_11_sva_1_39_16, and_dcpl_1118);
        attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_12_sva_1_39_16, and_dcpl_1121);
        attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_13_sva_1_39_16, and_dcpl_1124);
        attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_14_sva_1_39_16, and_dcpl_1127);
        attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_0_15_sva_1_39_16, and_dcpl_1130);
        attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0, and_dcpl_1084);
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_15_8 <= MUX_v_8_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 8)), APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8, and_dcpl_1088);
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_7 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(7)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7, and_dcpl_1088);
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_6 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(6)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6, and_dcpl_1088);
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_5 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(5)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5, and_dcpl_1088);
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_4 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(4)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4, and_dcpl_1088);
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_3 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(3)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3, and_dcpl_1088);
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_2 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(2)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2, and_dcpl_1088);
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_1 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(1)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1, and_dcpl_1088);
        attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_0 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(0)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0, and_dcpl_1088);
        attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_15_0, and_dcpl_1091);
        attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0,
            and_dcpl_1094);
        attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_15_0, and_dcpl_1097);
        attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_15_0, and_dcpl_1100);
        attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_15_0, and_dcpl_1103);
        attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0, and_dcpl_1106);
        attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_15_0, and_dcpl_1109);
        attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_15_0, and_dcpl_1112);
        attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_15_13 <= MUX_v_3_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 13)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd,
            and_dcpl_1115);
        attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0 <= MUX_v_13_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(12
            DOWNTO 0)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1,
            and_dcpl_1115);
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_15_8 <= MUX_v_8_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 8)), apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_15_8,
            and_dcpl_1118);
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_7 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(7)),
            apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_7, and_dcpl_1118);
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_6 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(6)),
            apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_6, and_dcpl_1118);
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_5 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(5)),
            apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_5, and_dcpl_1118);
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_4 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(4)),
            apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_4, and_dcpl_1118);
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_3 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(3)),
            apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_3, and_dcpl_1118);
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_2 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(2)),
            apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_2, and_dcpl_1118);
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_1 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(1)),
            apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_1, and_dcpl_1118);
        attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_0 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(0)),
            apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_0, and_dcpl_1118);
        attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0, and_dcpl_1121);
        attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_15_0, and_dcpl_1124);
        attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_15_0, and_dcpl_1127);
        attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0, and_dcpl_1130);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT(or_dcpl_1146
          OR and_dcpl_1055))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_v_proj_and_30_cse = '1' ) THEN
        attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16_mx0w5;
        attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0_mx0w6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva <= '0';
        GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva <= '0';
      ELSIF ( GEMM_3D_FLOAT_LOOP_3_1_and_44_cse = '1' ) THEN
        GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva <= MUX1HOT_s_1_4_2(APPLY_ROTARY_POS_EMB_LOOP_3_and_7_nl,
            GEMM_3D_FLOAT_LOOP_3_and_tmp_6_sva_mx0w1, GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva_mx0w3,
            (NOT QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1),
            STD_LOGIC_VECTOR'( and_dcpl_207 & and_dcpl_1152 & and_dcpl_222 & and_dcpl_1154));
        GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva <= MUX1HOT_s_1_4_2(APPLY_ROTARY_POS_EMB_LOOP_3_and_5_nl,
            GEMM_3D_FLOAT_LOOP_3_and_tmp_7_sva_mx0w1, GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva_mx0w3,
            QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1, STD_LOGIC_VECTOR'(
            and_dcpl_207 & and_dcpl_1152 & and_dcpl_222 & and_dcpl_1154));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_embed_3_0_3_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_3_0_2_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_3_0_1_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_3_0_0_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_q_embed_2_0_3_lpi_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_q_embed_and_cse = '1' ) THEN
        attention_2_1_16_16_4_4_q_embed_3_0_3_lpi_3 <= attention_2_1_16_16_4_4_q_embed_mux_14_cse;
        attention_2_1_16_16_4_4_q_embed_3_0_2_lpi_3 <= attention_2_1_16_16_4_4_q_embed_mux_13_cse;
        attention_2_1_16_16_4_4_q_embed_3_0_1_lpi_3 <= attention_2_1_16_16_4_4_q_embed_mux_11_cse;
        attention_2_1_16_16_4_4_q_embed_3_0_0_lpi_3 <= attention_2_1_16_16_4_4_q_embed_mux_9_cse;
        attention_2_1_16_16_4_4_q_embed_2_0_3_lpi_3 <= attention_2_1_16_16_4_4_q_embed_mux_7_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_q_embed_0_0_0_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT((NOT mux_2130_nl)
          AND and_dcpl_718))) = '1' ) THEN
        attention_2_1_16_16_4_4_q_embed_0_0_0_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
            attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1, or_dcpl_1025);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_k_embed_0_0_0_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT(mux_2131_nl
          AND (NOT (fsm_output(8))) AND and_dcpl_1145))) = '1' ) THEN
        attention_2_1_16_16_4_4_k_embed_0_0_0_sva_1 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_991)
          OR and_dcpl_346 OR attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c1
          OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_349 OR and_dcpl_351 OR and_dcpl_1162
          OR mux_tmp_2153 OR attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c9))
          = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            attention_2_1_16_16_4_4_q_embed_mux1h_40_nl, not_4510_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT(or_dcpl_996
          OR mux_2159_nl)) OR and_dcpl_346 OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_351
          OR mux_tmp_2176 OR attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx0c7))
          = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            attention_2_1_16_16_4_4_q_embed_mux1h_41_nl, not_4483_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT(or_dcpl_993
          OR mux_2182_nl)) OR and_dcpl_346 OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_351
          OR mux_tmp_2176 OR attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx0c7))
          = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            attention_2_1_16_16_4_4_q_embed_mux1h_42_nl, not_4482_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_990)
          OR and_dcpl_346 OR attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c1
          OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_349 OR and_dcpl_351 OR and_dcpl_1162
          OR mux_tmp_2153 OR attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c9))
          = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            attention_2_1_16_16_4_4_q_embed_mux1h_43_nl, not_4511_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_988)
          OR and_dcpl_346 OR mux_2198_nl OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_351
          OR mux_tmp_2176 OR attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx0c7)
          AND (and_dcpl_346 OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_351 OR mux_tmp_2176
          OR and_dcpl_352 OR attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx0c7))
          = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            attention_2_1_16_16_4_4_q_embed_mux1h_44_nl, not_4512_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_985)
          OR and_dcpl_346 OR mux_2204_nl OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_351
          OR mux_tmp_2176 OR attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx0c7)
          AND (and_dcpl_346 OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_351 OR mux_tmp_2176
          OR and_dcpl_352 OR attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx0c7))
          = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            attention_2_1_16_16_4_4_q_embed_mux1h_45_nl, not_4513_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_980)
          OR and_dcpl_346 OR mux_2210_nl OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_351
          OR mux_tmp_2176 OR attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx0c7)
          AND (and_dcpl_346 OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_351 OR mux_tmp_2176
          OR and_dcpl_352 OR attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx0c7))
          = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            attention_2_1_16_16_4_4_q_embed_mux1h_46_nl, not_4514_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_983)
          OR and_dcpl_346 OR attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c1
          OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_349 OR and_dcpl_351 OR and_dcpl_1162
          OR mux_tmp_2153 OR attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c9))
          = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            attention_2_1_16_16_4_4_q_embed_mux1h_47_nl, not_4515_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND ((NOT or_dcpl_987)
          OR and_dcpl_346 OR mux_2226_nl OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_351
          OR mux_tmp_2176 OR attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx0c7)
          AND (and_dcpl_346 OR and_dcpl_204 OR and_dcpl_348 OR and_dcpl_351 OR mux_tmp_2176
          OR and_dcpl_352 OR attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx0c7))
          = '1' ) THEN
        attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1 <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
            attention_2_1_16_16_4_4_q_embed_mux1h_48_nl, not_4516_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        TRANSPOSE_LAST_TWO_DIMS_LOOP_3_k_2_0_sva_1 <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT((NOT (fsm_output(0)))
          OR (NOT (fsm_output(1))) OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR
          (fsm_output(8)) OR or_dcpl_1134 OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")))))
          = '1' ) THEN
        TRANSPOSE_LAST_TWO_DIMS_LOOP_3_k_2_0_sva_1 <= z_out_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_attn_weights_and_cse = '1' ) THEN
        attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_35_nl,
            attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2_mx1, and_dcpl_193);
        attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_34_nl,
            attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2_mx1, and_dcpl_193);
        attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_33_nl,
            attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2_mx1, and_dcpl_193);
        attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_32_nl,
            attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2_mx1, and_dcpl_193);
        attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_31_nl,
            attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2_mx1, and_dcpl_193);
        attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_30_nl,
            attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2_mx1, and_dcpl_193);
        attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_29_nl,
            attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2_mx1, and_dcpl_193);
        attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_28_nl,
            attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2_mx1, and_dcpl_193);
        attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_27_nl,
            attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2_mx1, and_dcpl_193);
        attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_26_nl,
            attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2_mx1, and_dcpl_193);
        attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_25_nl,
            attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2_mx1, and_dcpl_193);
        attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_24_nl,
            attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2_mx1, and_dcpl_193);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        GEMM_3D_FLOAT_LOOP_3_and_tmp_sva <= '0';
        GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva <= '0';
        GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva <= '0';
        GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva <= '0';
        GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva <= '0';
        GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva <= '0';
        GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva <= '0';
        GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva <= '0';
      ELSIF ( GEMM_3D_FLOAT_LOOP_3_and_36_cse = '1' ) THEN
        GEMM_3D_FLOAT_LOOP_3_and_tmp_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_sva_mx0w0;
        GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva_mx0w0;
        GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva_mx0w0;
        GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva_mx0w0;
        GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva_mx0w0;
        GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva_mx0w0;
        GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva_mx0w0;
        GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_attn_weights_and_52_cse = '1' ) THEN
        attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1, and_dcpl_1199);
        attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1, and_dcpl_1199);
        attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1, and_dcpl_1199);
        attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1, and_dcpl_1199);
        attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1, and_dcpl_1199);
        attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1, and_dcpl_1199);
        attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1, and_dcpl_1199);
        attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1, and_dcpl_1199);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_3 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_attn_weights_and_48_cse = '1' ) THEN
        attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx1, and_dcpl_349);
        attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx1, and_dcpl_349);
        attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx1, and_dcpl_349);
        attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx1, and_dcpl_349);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_attn_weights_and_12_cse = '1' ) THEN
        attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_3,
            attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8_mx1, and_dcpl_377);
        attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1,
            attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9_mx1, and_dcpl_377);
        attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_3,
            attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8_mx1, and_dcpl_377);
        attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_3,
            attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8_mx1, and_dcpl_377);
        attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1,
            attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9_mx1, and_dcpl_377);
        attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_3,
            attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8_mx1, and_dcpl_377);
        attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_3,
            attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8_mx1, and_dcpl_377);
        attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1,
            attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9_mx1, and_dcpl_377);
        attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_3,
            attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8_mx1, and_dcpl_377);
        attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_3,
            attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8_mx1, and_dcpl_377);
        attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1,
            attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9_mx1, and_dcpl_377);
        attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_3,
            attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8_mx1, and_dcpl_377);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_4 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_5 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_4 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_4 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_5 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_4 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_4 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_5 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_4 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_4 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_5 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
        attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_4 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( attention_2_1_16_16_4_4_attn_weights_and_24_cse = '1' ) THEN
        attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx2, and_dcpl_351);
        attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_5 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx2, and_dcpl_351);
        attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx1, and_dcpl_351);
        attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx2, and_dcpl_351);
        attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_5 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx1, and_dcpl_351);
        attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx2, and_dcpl_351);
        attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx1, and_dcpl_351);
        attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_5 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx2, and_dcpl_351);
        attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx1, and_dcpl_351);
        attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx1, and_dcpl_351);
        attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_5 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx1, and_dcpl_351);
        attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8_mx1,
            attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx1, and_dcpl_351);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        softmax_1_4_3_sum_sva_1 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT(mux_2248_nl
          AND and_dcpl_295))) = '1' ) THEN
        softmax_1_4_3_sum_sva_1 <= softmax_1_4_3_sum_sva_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva <= '0';
        GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva <= '0';
        GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva <= '0';
        GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva <= '0';
      ELSIF ( GEMM_3D_FLOAT_LOOP_3_1_and_46_cse = '1' ) THEN
        GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva <= GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva_mx0w0;
        GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva <= GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva_mx0w0;
        GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva <= GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva_mx0w0;
        GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva <= GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_abs_4_qr_35_0_lpi_1_dfm_35 <= '0';
        attention_abs_4_qr_35_0_lpi_1_dfm_34_0 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000");
      ELSIF ( attention_abs_4_qelse_and_ssc = '1' ) THEN
        attention_abs_4_qr_35_0_lpi_1_dfm_35 <= (attention_abs_qr_35_0_lpi_1_dfm_mx0w0(35))
            AND (NOT attention_abs_4_qr_35_0_lpi_1_dfm_mx0c1);
        attention_abs_4_qr_35_0_lpi_1_dfm_34_0 <= MUX_v_35_2_2((attention_abs_qr_35_0_lpi_1_dfm_mx0w0(34
            DOWNTO 0)), (operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1(34
            DOWNTO 0)), attention_abs_4_qr_35_0_lpi_1_dfm_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        compute_sqrt_1_guess_sva_34 <= '0';
        compute_sqrt_1_guess_sva_33_0 <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000");
      ELSIF ( compute_sqrt_1_guess_and_ssc = '1' ) THEN
        compute_sqrt_1_guess_sva_34 <= MUX_s_1_2_2(attention_abs_qr_35_0_lpi_1_dfm_mx1_35,
            (compute_sqrt_1_for_acc_1_itm_40_1_1(34)), and_dcpl_292);
        compute_sqrt_1_guess_sva_33_0 <= MUX_v_34_2_2(attention_abs_qr_35_0_lpi_1_dfm_mx1_34_1,
            (compute_sqrt_1_for_acc_1_itm_40_1_1(33 DOWNTO 0)), and_dcpl_292);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_38_0 <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND and_dcpl_548)
          = '1' ) THEN
        QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_38_0 <= QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_dfm_1_38_0_mx0w1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_cse = '1' ) THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
        attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_8_cse = '1' ) THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
        attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_16_cse = '1' ) THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
        attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_24_cse = '1' ) THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
        attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_32_cse = '1' ) THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
        attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_40_cse = '1' ) THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
        attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_48_cse = '1' ) THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
        attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_56_cse = '1' ) THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
        attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_64_cse = '1' ) THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
        attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_72_cse = '1' ) THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
        attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_80_cse = '1' ) THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
        attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_88_cse = '1' ) THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
        attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_96_cse = '1' ) THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
        attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_7 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_104_cse = '1' )
          THEN
        reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
        attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva <= STD_LOGIC_VECTOR'(
            "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT(or_tmp_833
          OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR or_dcpl_1109
          OR nand_253_cse))) = '1' ) THEN
        RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva <= z_out_13_71_28(43
            DOWNTO 4);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT and_dcpl_414))
          = '1' ) THEN
        QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva <= LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
            DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_7 <= '0';
        attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3 <= '0';
      ELSIF ( attention_2_1_16_16_4_4_quantized_final_output_and_112_cse = '1' )
          THEN
        attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_7 <= NOT((NOT QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1)
            OR QUANTIZE_ACTIVATION_LOOP_3_1_nand_seb_1);
        attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3 <= NOT(QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1
            OR QUANTIZE_ACTIVATION_LOOP_3_1_nand_seb_1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_0_15_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_0_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_14_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_1_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_13_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_2_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_12_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_3_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_11_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_4_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_10_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_5_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_9_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_6_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_8_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
        output_0_7_sva_1_39_16 <= STD_LOGIC_VECTOR'( "000000000000000000000000");
      ELSIF ( output_and_16_cse = '1' ) THEN
        output_0_15_sva_1_39_16 <= output_0_15_lpi_4_39_16_mx1;
        output_0_0_sva_1_39_16 <= output_0_0_lpi_4_39_16_mx1;
        output_0_14_sva_1_39_16 <= output_0_14_lpi_4_39_16_mx1;
        output_0_1_sva_1_39_16 <= output_0_1_lpi_4_39_16_mx1;
        output_0_13_sva_1_39_16 <= output_0_13_lpi_4_39_16_mx1;
        output_0_2_sva_1_39_16 <= output_0_2_lpi_4_39_16_mx1;
        output_0_12_sva_1_39_16 <= output_0_12_lpi_4_39_16_mx1;
        output_0_3_sva_1_39_16 <= output_0_3_lpi_4_39_16_mx1;
        output_0_11_sva_1_39_16 <= output_0_11_lpi_4_39_16_mx1;
        output_0_4_sva_1_39_16 <= output_0_4_lpi_4_39_16_mx1;
        output_0_10_sva_1_39_16 <= output_0_10_lpi_4_39_16_mx1;
        output_0_5_sva_1_39_16 <= output_0_5_lpi_4_39_16_mx1;
        output_0_9_sva_1_39_16 <= output_0_9_lpi_4_39_16_mx1;
        output_0_6_sva_1_39_16 <= output_0_6_lpi_4_39_16_mx1;
        output_0_8_sva_1_39_16 <= output_0_8_lpi_4_39_16_mx1;
        output_0_7_sva_1_39_16 <= output_0_7_lpi_4_39_16_mx1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        LINEAR_FORWARD_NO_MUL_LOOP_2_3_mul_mut <= STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000000000000000000000000");
      ELSIF ( (attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 AND (NOT(or_dcpl_961
          OR or_dcpl_1134 OR or_1984_cse))) = '1' ) THEN
        LINEAR_FORWARD_NO_MUL_LOOP_2_3_mul_mut <= z_out_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_0_0_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_1_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_2_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_3_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_4_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_5_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_6_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_7_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_8_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_9_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_10_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_11_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_12_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_13_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_14_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_15_sva_2_29_16 <= STD_LOGIC_VECTOR'( "00000000000000");
        output_0_0_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_1_sva_2_15_8 <= STD_LOGIC_VECTOR'( "00000000");
        output_0_1_sva_2_7 <= '0';
        output_0_1_sva_2_6 <= '0';
        output_0_1_sva_2_5 <= '0';
        output_0_1_sva_2_4 <= '0';
        output_0_1_sva_2_3 <= '0';
        output_0_1_sva_2_2 <= '0';
        output_0_1_sva_2_1 <= '0';
        output_0_1_sva_2_0 <= '0';
        output_0_2_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_3_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_4_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_5_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_6_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_7_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_8_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_9_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_10_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_11_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_12_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_13_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_14_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
        output_0_15_sva_2_15_0 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( output_and_64_cse = '1' ) THEN
        output_0_0_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_0_sva_1_39_16(13 DOWNTO 0)), output_and_35_nl);
        output_0_1_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_1_sva_1_39_16(13 DOWNTO 0)), output_and_39_nl);
        output_0_2_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_2_sva_1_39_16(13 DOWNTO 0)), output_and_43_nl);
        output_0_3_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_3_sva_1_39_16(13 DOWNTO 0)), output_and_47_nl);
        output_0_4_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_4_sva_1_39_16(13 DOWNTO 0)), output_and_51_nl);
        output_0_5_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_5_sva_1_39_16(13 DOWNTO 0)), output_and_55_nl);
        output_0_6_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_6_sva_1_39_16(13 DOWNTO 0)), output_and_59_nl);
        output_0_7_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_7_sva_1_39_16(13 DOWNTO 0)), output_and_63_nl);
        output_0_8_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_8_sva_1_39_16(13 DOWNTO 0)), output_and_61_nl);
        output_0_9_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_9_sva_1_39_16(13 DOWNTO 0)), output_and_57_nl);
        output_0_10_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_10_sva_1_39_16(13 DOWNTO 0)), output_and_53_nl);
        output_0_11_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_11_sva_1_39_16(13 DOWNTO 0)), output_and_49_nl);
        output_0_12_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_12_sva_1_39_16(13 DOWNTO 0)), output_and_45_nl);
        output_0_13_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_13_sva_1_39_16(13 DOWNTO 0)), output_and_41_nl);
        output_0_14_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_14_sva_1_39_16(13 DOWNTO 0)), output_and_37_nl);
        output_0_15_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(29
            DOWNTO 16)), (output_0_15_sva_1_39_16(13 DOWNTO 0)), output_and_33_nl);
        output_0_0_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0, or_dcpl_1155);
        output_0_1_sva_2_15_8 <= MUX_v_8_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 8)), APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8, or_dcpl_1158);
        output_0_1_sva_2_7 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(7)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7, or_dcpl_1158);
        output_0_1_sva_2_6 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(6)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6, or_dcpl_1158);
        output_0_1_sva_2_5 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(5)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5, or_dcpl_1158);
        output_0_1_sva_2_4 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(4)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4, or_dcpl_1158);
        output_0_1_sva_2_3 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(3)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3, or_dcpl_1158);
        output_0_1_sva_2_2 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(2)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2, or_dcpl_1158);
        output_0_1_sva_2_1 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(1)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1, or_dcpl_1158);
        output_0_1_sva_2_0 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(0)),
            APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0, or_dcpl_1158);
        output_0_2_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0,
            or_dcpl_1160);
        output_0_3_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0,
            or_dcpl_1162);
        output_0_4_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0, or_dcpl_1165);
        output_0_5_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0, or_dcpl_1167);
        output_0_6_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0, or_dcpl_1169);
        output_0_7_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0, or_dcpl_1141);
        output_0_8_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0, or_dcpl_1170);
        output_0_9_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0, or_dcpl_1168);
        output_0_10_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0, or_dcpl_1166);
        output_0_11_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0, or_dcpl_1164);
        output_0_12_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0, or_dcpl_1161);
        output_0_13_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0, or_dcpl_1159);
        output_0_14_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0, or_dcpl_1156);
        output_0_15_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
            DOWNTO 0)), attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0, or_dcpl_1152);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd <= '0';
        reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 <= '0';
      ELSIF ( GEMM_3D_FLOAT_LOOP_4_l_and_ssc = '1' ) THEN
        reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd <= GEMM_3D_FLOAT_LOOP_4_l_mux1h_6_nl
            AND (NOT GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c2);
        reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 <= GEMM_3D_FLOAT_LOOP_4_l_mux1h_8_nl
            AND (NOT GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c2);
      END IF;
    END IF;
  END PROCESS;
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_nl <= MUX1HOT_v_8_4_2((drf_output_sdt_2_sva_15_0_mx0w0(15
      DOWNTO 8)), reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd, (drf_output_sdt_3_sva_15_0_mx0w3(15
      DOWNTO 8)), LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8, STD_LOGIC_VECTOR'(
      and_dcpl_257 & and_dcpl_260 & and_dcpl_265 & and_dcpl_268));
  not_4947_nl <= NOT or_dcpl_1048;
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_1_nl <= MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0(7)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7, (drf_output_sdt_3_sva_15_0_mx0w3(7)),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd, STD_LOGIC_VECTOR'( and_dcpl_257
      & and_dcpl_260 & and_dcpl_265 & and_dcpl_268));
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_2_nl <= MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0(6)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6, (drf_output_sdt_3_sva_15_0_mx0w3(6)),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1, STD_LOGIC_VECTOR'( and_dcpl_257
      & and_dcpl_260 & and_dcpl_265 & and_dcpl_268));
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_3_nl <= MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0(5)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5, (drf_output_sdt_3_sva_15_0_mx0w3(5)),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2, STD_LOGIC_VECTOR'( and_dcpl_257
      & and_dcpl_260 & and_dcpl_265 & and_dcpl_268));
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_4_nl <= MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0(4)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4, (drf_output_sdt_3_sva_15_0_mx0w3(4)),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3, STD_LOGIC_VECTOR'( and_dcpl_257
      & and_dcpl_260 & and_dcpl_265 & and_dcpl_268));
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_5_nl <= MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0(3)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3, (drf_output_sdt_3_sva_15_0_mx0w3(3)),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4, STD_LOGIC_VECTOR'( and_dcpl_257
      & and_dcpl_260 & and_dcpl_265 & and_dcpl_268));
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_6_nl <= MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0(2)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2, (drf_output_sdt_3_sva_15_0_mx0w3(2)),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5, STD_LOGIC_VECTOR'( and_dcpl_257
      & and_dcpl_260 & and_dcpl_265 & and_dcpl_268));
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_7_nl <= MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0(1)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1, (drf_output_sdt_3_sva_15_0_mx0w3(1)),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6, STD_LOGIC_VECTOR'( and_dcpl_257
      & and_dcpl_260 & and_dcpl_265 & and_dcpl_268));
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_8_nl <= MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0(0)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0, (drf_output_sdt_3_sva_15_0_mx0w3(0)),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7, STD_LOGIC_VECTOR'( and_dcpl_257
      & and_dcpl_260 & and_dcpl_265 & and_dcpl_268));
  rms_norm_16_mux1h_nl <= MUX1HOT_s_1_5_2(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4,
      (compute_sqrt_for_acc_1_itm_40_1_1(39)), attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_39,
      reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd, (compute_sqrt_1_for_acc_1_itm_40_1_1(39)),
      STD_LOGIC_VECTOR'( and_321_ssc & and_dcpl_290 & and_dcpl_276 & and_dcpl_278
      & and_dcpl_292));
  rms_norm_16_mux1h_9_nl <= MUX1HOT_v_4_5_2(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0,
      (compute_sqrt_for_acc_1_itm_40_1_1(38 DOWNTO 35)), (attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_38_0(38
      DOWNTO 35)), (reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(38 DOWNTO 35)), (compute_sqrt_1_for_acc_1_itm_40_1_1(38
      DOWNTO 35)), STD_LOGIC_VECTOR'( and_321_ssc & and_dcpl_290 & and_dcpl_276 &
      and_dcpl_278 & and_dcpl_292));
  operator_40_24_true_AC_TRN_AC_WRAP_1_not_1_nl <= NOT mux_851_ssc;
  SOFTMAX_LOOP_5_mux_24_nl <= MUX_s_1_2_2((SOFTMAX_LOOP_5_mux_12_psp_mx0w0(39)),
      reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd, and_329_ssc);
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_mux1h_2_nl <= MUX1HOT_v_24_4_2(LINEAR_FORWARD_NO_MUL_LOOP_2_2_conc_1_mut_71_48_mx0w0,
      for_for_strm_in_tmp_sva_25_2, LINEAR_FORWARD_NO_MUL_LOOP_2_3_conc_1_mut_71_48_mx0w3,
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48, STD_LOGIC_VECTOR'( and_dcpl_257
      & and_dcpl_260 & and_dcpl_265 & and_dcpl_268));
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_not_nl <= NOT or_dcpl_1048;
  mux_862_nl <= MUX_s_1_2_2((NOT mux_tmp_787), or_1732_cse, for_for_and_tmp);
  rms_norm_16_mux1h_10_nl <= MUX1HOT_s_1_4_2((compute_sqrt_for_acc_1_itm_40_1_1(0)),
      (reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(0)), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2(0)),
      (LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut(0)), STD_LOGIC_VECTOR'( and_dcpl_290
      & and_343_itm & and_dcpl_257 & and_dcpl_260));
  rms_norm_16_mux1h_6_nl <= MUX1HOT_v_24_3_2(LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48_mx0w2,
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48, APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16,
      STD_LOGIC_VECTOR'( and_dcpl_257 & and_dcpl_260 & and_dcpl_310));
  rms_norm_16_not_nl <= NOT rms_norm_16_div_cmp_a_mx0c0;
  rms_norm_16_mux1h_7_nl <= MUX1HOT_v_8_3_2((z_out_1(15 DOWNTO 8)), LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd, STD_LOGIC_VECTOR'( and_dcpl_257
      & and_dcpl_260 & and_dcpl_310));
  rms_norm_16_not_1_nl <= NOT rms_norm_16_div_cmp_a_mx0c0;
  rms_norm_16_mux1h_11_nl <= MUX1HOT_s_1_3_2((z_out_1(7)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7, STD_LOGIC_VECTOR'(
      and_dcpl_257 & and_dcpl_260 & and_dcpl_310));
  rms_norm_16_mux1h_13_nl <= MUX1HOT_s_1_3_2((z_out_1(6)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6, STD_LOGIC_VECTOR'(
      and_dcpl_257 & and_dcpl_260 & and_dcpl_310));
  rms_norm_16_mux1h_14_nl <= MUX1HOT_s_1_3_2((z_out_1(5)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5, STD_LOGIC_VECTOR'(
      and_dcpl_257 & and_dcpl_260 & and_dcpl_310));
  rms_norm_16_mux1h_15_nl <= MUX1HOT_s_1_3_2((z_out_1(4)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4, STD_LOGIC_VECTOR'(
      and_dcpl_257 & and_dcpl_260 & and_dcpl_310));
  rms_norm_16_mux1h_16_nl <= MUX1HOT_s_1_3_2((z_out_1(3)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3, STD_LOGIC_VECTOR'(
      and_dcpl_257 & and_dcpl_260 & and_dcpl_310));
  rms_norm_16_mux1h_17_nl <= MUX1HOT_s_1_3_2((z_out_1(2)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2, STD_LOGIC_VECTOR'(
      and_dcpl_257 & and_dcpl_260 & and_dcpl_310));
  rms_norm_16_mux1h_18_nl <= MUX1HOT_s_1_3_2((z_out_1(1)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1, STD_LOGIC_VECTOR'(
      and_dcpl_257 & and_dcpl_260 & and_dcpl_310));
  rms_norm_16_mux1h_19_nl <= MUX1HOT_s_1_3_2((z_out_1(0)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0, STD_LOGIC_VECTOR'(
      and_dcpl_257 & and_dcpl_260 & and_dcpl_310));
  INIT_2D_MEM_LOOP_2_mux_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_633_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_nl <= INIT_2D_MEM_LOOP_2_mux_nl AND (NOT
      or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_10_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_633_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_38_nl <= INIT_2D_MEM_LOOP_2_mux_10_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_11_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_633_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_39_nl <= INIT_2D_MEM_LOOP_2_mux_11_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_12_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_633_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_40_nl <= INIT_2D_MEM_LOOP_2_mux_12_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_13_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_633_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_41_nl <= INIT_2D_MEM_LOOP_2_mux_13_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_14_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_633_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_42_nl <= INIT_2D_MEM_LOOP_2_mux_14_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_15_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_633_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_43_nl <= INIT_2D_MEM_LOOP_2_mux_15_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_16_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_633_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_44_nl <= INIT_2D_MEM_LOOP_2_mux_16_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_1_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_654_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_1_nl <= INIT_2D_MEM_LOOP_2_mux_1_nl AND
      (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_17_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_654_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_24_nl <= INIT_2D_MEM_LOOP_2_mux_17_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_18_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_654_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_nl <= INIT_2D_MEM_LOOP_2_mux_18_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_19_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_654_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_26_nl <= INIT_2D_MEM_LOOP_2_mux_19_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_20_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_654_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_27_nl <= INIT_2D_MEM_LOOP_2_mux_20_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_21_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_654_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_28_nl <= INIT_2D_MEM_LOOP_2_mux_21_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_22_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_654_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_29_nl <= INIT_2D_MEM_LOOP_2_mux_22_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_23_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_654_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_30_nl <= INIT_2D_MEM_LOOP_2_mux_23_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_2_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_648_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_2_nl <= INIT_2D_MEM_LOOP_2_mux_2_nl AND
      (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_24_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_648_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_10_nl <= INIT_2D_MEM_LOOP_2_mux_24_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_25_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_648_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_11_nl <= INIT_2D_MEM_LOOP_2_mux_25_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_26_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_648_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_12_nl <= INIT_2D_MEM_LOOP_2_mux_26_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_27_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_648_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_13_nl <= INIT_2D_MEM_LOOP_2_mux_27_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_28_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_648_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_14_nl <= INIT_2D_MEM_LOOP_2_mux_28_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_29_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_648_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_15_nl <= INIT_2D_MEM_LOOP_2_mux_29_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_30_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_648_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_16_nl <= INIT_2D_MEM_LOOP_2_mux_30_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_3_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_642_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_3_nl <= INIT_2D_MEM_LOOP_2_mux_3_nl AND
      (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_31_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_642_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_17_nl <= INIT_2D_MEM_LOOP_2_mux_31_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_32_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_642_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_18_nl <= INIT_2D_MEM_LOOP_2_mux_32_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_33_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_642_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_19_nl <= INIT_2D_MEM_LOOP_2_mux_33_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_34_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_642_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_20_nl <= INIT_2D_MEM_LOOP_2_mux_34_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_35_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_642_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_21_nl <= INIT_2D_MEM_LOOP_2_mux_35_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_36_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_642_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_22_nl <= INIT_2D_MEM_LOOP_2_mux_36_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_37_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_642_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_23_nl <= INIT_2D_MEM_LOOP_2_mux_37_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_4_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_636_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_4_nl <= INIT_2D_MEM_LOOP_2_mux_4_nl AND
      (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_38_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_636_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_31_nl <= INIT_2D_MEM_LOOP_2_mux_38_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_39_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_636_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_32_nl <= INIT_2D_MEM_LOOP_2_mux_39_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_40_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_636_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_33_nl <= INIT_2D_MEM_LOOP_2_mux_40_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_41_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_636_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_34_nl <= INIT_2D_MEM_LOOP_2_mux_41_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_42_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_636_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_35_nl <= INIT_2D_MEM_LOOP_2_mux_42_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_43_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_636_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_36_nl <= INIT_2D_MEM_LOOP_2_mux_43_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_44_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_636_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_37_nl <= INIT_2D_MEM_LOOP_2_mux_44_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_5_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_629_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_5_nl <= INIT_2D_MEM_LOOP_2_mux_5_nl AND
      (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_45_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_629_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_45_nl <= INIT_2D_MEM_LOOP_2_mux_45_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_46_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_629_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_46_nl <= INIT_2D_MEM_LOOP_2_mux_46_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_47_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_629_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_47_nl <= INIT_2D_MEM_LOOP_2_mux_47_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_48_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_629_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_48_nl <= INIT_2D_MEM_LOOP_2_mux_48_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_49_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_629_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_49_nl <= INIT_2D_MEM_LOOP_2_mux_49_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_50_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_629_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_50_nl <= INIT_2D_MEM_LOOP_2_mux_50_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_51_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_629_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_51_nl <= INIT_2D_MEM_LOOP_2_mux_51_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_6_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_639_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_6_nl <= INIT_2D_MEM_LOOP_2_mux_6_nl AND
      (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_52_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_639_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_52_nl <= INIT_2D_MEM_LOOP_2_mux_52_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_53_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_639_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_53_nl <= INIT_2D_MEM_LOOP_2_mux_53_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_54_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_639_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_54_nl <= INIT_2D_MEM_LOOP_2_mux_54_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_55_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_639_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_55_nl <= INIT_2D_MEM_LOOP_2_mux_55_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_56_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_639_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_56_nl <= INIT_2D_MEM_LOOP_2_mux_56_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_57_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_639_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_57_nl <= INIT_2D_MEM_LOOP_2_mux_57_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_58_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_639_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_58_nl <= INIT_2D_MEM_LOOP_2_mux_58_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_7_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_645_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_7_nl <= INIT_2D_MEM_LOOP_2_mux_7_nl AND
      (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_59_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_645_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_59_nl <= INIT_2D_MEM_LOOP_2_mux_59_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_60_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_645_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_60_nl <= INIT_2D_MEM_LOOP_2_mux_60_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_61_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_645_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_61_nl <= INIT_2D_MEM_LOOP_2_mux_61_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_62_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_645_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_62_nl <= INIT_2D_MEM_LOOP_2_mux_62_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_63_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_645_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_63_nl <= INIT_2D_MEM_LOOP_2_mux_63_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_64_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_645_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_64_nl <= INIT_2D_MEM_LOOP_2_mux_64_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_65_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_645_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_65_nl <= INIT_2D_MEM_LOOP_2_mux_65_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_8_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_651_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_8_nl <= INIT_2D_MEM_LOOP_2_mux_8_nl AND
      (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_66_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_651_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_66_nl <= INIT_2D_MEM_LOOP_2_mux_66_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_67_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_651_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_67_nl <= INIT_2D_MEM_LOOP_2_mux_67_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_68_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_651_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_68_nl <= INIT_2D_MEM_LOOP_2_mux_68_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_69_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_651_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_69_nl <= INIT_2D_MEM_LOOP_2_mux_69_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_70_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_651_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_70_nl <= INIT_2D_MEM_LOOP_2_mux_70_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_71_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_651_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_71_nl <= INIT_2D_MEM_LOOP_2_mux_71_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_72_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_651_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_72_nl <= INIT_2D_MEM_LOOP_2_mux_72_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_9_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_657_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_9_nl <= INIT_2D_MEM_LOOP_2_mux_9_nl AND
      (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_73_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_657_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_73_nl <= INIT_2D_MEM_LOOP_2_mux_73_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_74_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_657_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_74_nl <= INIT_2D_MEM_LOOP_2_mux_74_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_75_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_657_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_75_nl <= INIT_2D_MEM_LOOP_2_mux_75_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_76_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_657_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_76_nl <= INIT_2D_MEM_LOOP_2_mux_76_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_77_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_657_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_77_nl <= INIT_2D_MEM_LOOP_2_mux_77_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_78_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_657_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_78_nl <= INIT_2D_MEM_LOOP_2_mux_78_nl
      AND (NOT or_dcpl_1104);
  INIT_2D_MEM_LOOP_2_mux_79_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_657_itm);
  INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_79_nl <= INIT_2D_MEM_LOOP_2_mux_79_nl
      AND (NOT or_dcpl_1104);
  and_779_nl <= and_dcpl_732 AND and_dcpl_730;
  and_1653_nl <= (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd) AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      AND CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2=STD_LOGIC_VECTOR'("11"));
  mux_1556_nl <= MUX_s_1_2_2(mux_1555_cse, mux_1553_cse, and_1653_nl);
  mux_1558_nl <= MUX_s_1_2_2(mux_1557_cse, mux_1556_nl, fsm_output(0));
  mux_1560_nl <= MUX_s_1_2_2(mux_1559_cse, mux_1558_nl, and_1773_cse);
  mux_1561_nl <= MUX_s_1_2_2(mux_1560_nl, mux_1546_cse, fsm_output(7));
  and_783_nl <= and_dcpl_736 AND and_dcpl_730;
  and_790_nl <= and_dcpl_743 AND and_dcpl_740 AND and_dcpl_728;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_5_nl <= MUX1HOT_v_16_5_2(z_out_1, attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0,
      (rms_norm_16_div_cmp_z_oreg(15 DOWNTO 0)), output_0_7_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      STD_LOGIC_VECTOR'( and_779_nl & (NOT mux_1561_nl) & and_783_nl & and_dcpl_739
      & and_790_nl));
  not_4472_nl <= NOT and_dcpl_619;
  and_943_nl <= and_dcpl_732 AND and_dcpl_842;
  nor_466_nl <= NOT((NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd) OR
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("10")));
  mux_1655_nl <= MUX_s_1_2_2(mux_1555_cse, mux_1553_cse, nor_466_nl);
  mux_1657_nl <= MUX_s_1_2_2(mux_1557_cse, mux_1655_nl, fsm_output(0));
  mux_1659_nl <= MUX_s_1_2_2(mux_1559_cse, mux_1657_nl, and_1773_cse);
  mux_1660_nl <= MUX_s_1_2_2(mux_1659_nl, mux_1645_cse, fsm_output(7));
  attention_2_1_16_16_4_4_k_proj_re_nand_nl <= NOT(mux_1660_nl AND (NOT(or_dcpl_1010
      AND and_dcpl_207)));
  attention_2_1_16_16_4_4_k_proj_re_and_81_nl <= (NOT or_dcpl_1010) AND and_dcpl_207;
  and_945_nl <= and_dcpl_743 AND and_dcpl_551 AND and_dcpl_841;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_30_nl <= MUX1HOT_v_16_7_2(z_out_1, attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0,
      (rms_norm_16_div_cmp_z_oreg(15 DOWNTO 0)), RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_15_0, output_0_10_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      STD_LOGIC_VECTOR'( and_943_nl & attention_2_1_16_16_4_4_k_proj_re_nand_nl &
      and_dcpl_843 & attention_2_1_16_16_4_4_k_proj_re_and_81_nl & and_dcpl_847 &
      and_dcpl_739 & and_945_nl));
  not_4469_nl <= NOT and_dcpl_619;
  and_946_nl <= and_dcpl_732 AND and_dcpl_855;
  and_1684_nl <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd AND (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1)
      AND CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2=STD_LOGIC_VECTOR'("11"));
  mux_1671_nl <= MUX_s_1_2_2(mux_1555_cse, mux_1553_cse, and_1684_nl);
  mux_1673_nl <= MUX_s_1_2_2(mux_1557_cse, mux_1671_nl, fsm_output(0));
  mux_1675_nl <= MUX_s_1_2_2(mux_1559_cse, mux_1673_nl, and_1773_cse);
  mux_1676_nl <= MUX_s_1_2_2(mux_1675_nl, mux_1645_cse, fsm_output(7));
  attention_2_1_16_16_4_4_k_proj_re_nand_2_nl <= NOT(mux_1676_nl AND (NOT(or_dcpl_1012
      AND and_dcpl_207)));
  attention_2_1_16_16_4_4_k_proj_re_and_83_nl <= (NOT or_dcpl_1012) AND and_dcpl_207;
  and_948_nl <= and_dcpl_743 AND and_dcpl_551 AND and_dcpl_854;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_32_nl <= MUX1HOT_v_16_7_2(z_out_1, attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0,
      (rms_norm_16_div_cmp_z_oreg(15 DOWNTO 0)), RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_15_0, output_0_11_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      STD_LOGIC_VECTOR'( and_946_nl & attention_2_1_16_16_4_4_k_proj_re_nand_2_nl
      & and_dcpl_856 & attention_2_1_16_16_4_4_k_proj_re_and_83_nl & and_dcpl_847
      & and_dcpl_739 & and_948_nl));
  not_4468_nl <= NOT and_dcpl_619;
  and_949_nl <= and_dcpl_732 AND and_dcpl_859;
  or_2589_nl <= (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd) OR (NOT
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1) OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("00"));
  mux_1687_nl <= MUX_s_1_2_2(mux_1553_cse, mux_1555_cse, or_2589_nl);
  mux_1689_nl <= MUX_s_1_2_2(mux_1557_cse, mux_1687_nl, fsm_output(0));
  mux_1691_nl <= MUX_s_1_2_2(mux_1559_cse, mux_1689_nl, and_1773_cse);
  mux_1692_nl <= MUX_s_1_2_2(mux_1691_nl, mux_1645_cse, fsm_output(7));
  attention_2_1_16_16_4_4_k_proj_re_nand_4_nl <= NOT(mux_1692_nl AND (NOT(or_dcpl_1014
      AND and_dcpl_207)));
  attention_2_1_16_16_4_4_k_proj_re_and_85_nl <= (NOT or_dcpl_1014) AND and_dcpl_207;
  and_951_nl <= and_dcpl_743 AND and_dcpl_740 AND and_dcpl_818;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_34_nl <= MUX1HOT_v_16_7_2(z_out_1, attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0,
      (rms_norm_16_div_cmp_z_oreg(15 DOWNTO 0)), RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_15_0, output_0_12_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      STD_LOGIC_VECTOR'( and_949_nl & attention_2_1_16_16_4_4_k_proj_re_nand_4_nl
      & and_dcpl_860 & attention_2_1_16_16_4_4_k_proj_re_and_85_nl & and_dcpl_847
      & and_dcpl_739 & and_951_nl));
  not_4467_nl <= NOT and_dcpl_619;
  and_952_nl <= and_dcpl_732 AND and_dcpl_863;
  nand_367_nl <= NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      AND CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2=STD_LOGIC_VECTOR'("01")));
  mux_1703_nl <= MUX_s_1_2_2(mux_1553_cse, mux_1555_cse, nand_367_nl);
  mux_1705_nl <= MUX_s_1_2_2(mux_1557_cse, mux_1703_nl, fsm_output(0));
  mux_1707_nl <= MUX_s_1_2_2(mux_1559_cse, mux_1705_nl, and_1773_cse);
  mux_1708_nl <= MUX_s_1_2_2(mux_1707_nl, mux_1645_cse, fsm_output(7));
  attention_2_1_16_16_4_4_k_proj_re_nand_6_nl <= NOT(mux_1708_nl AND (NOT(or_dcpl_1016
      AND and_dcpl_207)));
  attention_2_1_16_16_4_4_k_proj_re_and_87_nl <= (NOT or_dcpl_1016) AND and_dcpl_207;
  and_954_nl <= and_dcpl_743 AND and_dcpl_740 AND and_dcpl_830;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_36_nl <= MUX1HOT_v_16_7_2(z_out_1, attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0,
      (rms_norm_16_div_cmp_z_oreg(15 DOWNTO 0)), RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_15_0, output_0_13_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      STD_LOGIC_VECTOR'( and_952_nl & attention_2_1_16_16_4_4_k_proj_re_nand_6_nl
      & and_dcpl_864 & attention_2_1_16_16_4_4_k_proj_re_and_87_nl & and_dcpl_847
      & and_dcpl_739 & and_954_nl));
  not_4466_nl <= NOT and_dcpl_619;
  and_955_nl <= and_dcpl_732 AND and_dcpl_871;
  and_1697_nl <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      AND CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2=STD_LOGIC_VECTOR'("10"));
  mux_1719_nl <= MUX_s_1_2_2(mux_1555_cse, mux_1553_cse, and_1697_nl);
  mux_1721_nl <= MUX_s_1_2_2(mux_1557_cse, mux_1719_nl, fsm_output(0));
  mux_1723_nl <= MUX_s_1_2_2(mux_1559_cse, mux_1721_nl, and_1773_cse);
  mux_1724_nl <= MUX_s_1_2_2(mux_1723_nl, mux_1645_cse, fsm_output(7));
  attention_2_1_16_16_4_4_k_proj_re_nand_8_nl <= NOT(mux_1724_nl AND (NOT(or_dcpl_1018
      AND and_dcpl_207)));
  attention_2_1_16_16_4_4_k_proj_re_and_89_nl <= (NOT or_dcpl_1018) AND and_dcpl_207;
  and_957_nl <= and_dcpl_743 AND and_dcpl_740 AND and_dcpl_841;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_38_nl <= MUX1HOT_v_16_7_2(z_out_1, attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0,
      (rms_norm_16_div_cmp_z_oreg(15 DOWNTO 0)), RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_15_0, output_0_14_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      STD_LOGIC_VECTOR'( and_955_nl & attention_2_1_16_16_4_4_k_proj_re_nand_8_nl
      & and_dcpl_872 & attention_2_1_16_16_4_4_k_proj_re_and_89_nl & and_dcpl_847
      & and_dcpl_739 & and_957_nl));
  not_4465_nl <= NOT and_dcpl_619;
  and_960_nl <= and_dcpl_732 AND and_dcpl_850;
  or_2611_nl <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd OR (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1)
      OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("00"));
  mux_1738_nl <= MUX_s_1_2_2(mux_1553_cse, mux_1555_cse, or_2611_nl);
  mux_1740_nl <= MUX_s_1_2_2(mux_1557_cse, mux_1738_nl, fsm_output(0));
  mux_1742_nl <= MUX_s_1_2_2(mux_1559_cse, mux_1740_nl, and_1773_cse);
  mux_1743_nl <= MUX_s_1_2_2(mux_1742_nl, mux_1546_cse, fsm_output(7));
  and_962_nl <= and_dcpl_743 AND and_dcpl_740 AND and_dcpl_550;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_42_nl <= MUX1HOT_v_16_5_2(z_out_1, attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0,
      (rms_norm_16_div_cmp_z_oreg(15 DOWNTO 0)), output_0_4_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      STD_LOGIC_VECTOR'( and_960_nl & (NOT mux_1743_nl) & and_dcpl_851 & and_dcpl_739
      & and_962_nl));
  not_4463_nl <= NOT and_dcpl_619;
  and_963_nl <= and_dcpl_732 AND and_dcpl_836;
  or_2617_nl <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd OR (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1)
      OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("01"));
  mux_1754_nl <= MUX_s_1_2_2(mux_1553_cse, mux_1555_cse, or_2617_nl);
  mux_1756_nl <= MUX_s_1_2_2(mux_1557_cse, mux_1754_nl, fsm_output(0));
  mux_1758_nl <= MUX_s_1_2_2(mux_1559_cse, mux_1756_nl, and_1773_cse);
  mux_1759_nl <= MUX_s_1_2_2(mux_1758_nl, mux_1546_cse, fsm_output(7));
  and_965_nl <= and_dcpl_743 AND and_dcpl_740 AND and_dcpl_835;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_44_nl <= MUX1HOT_v_16_5_2(z_out_1, attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0,
      (rms_norm_16_div_cmp_z_oreg(15 DOWNTO 0)), output_0_5_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      STD_LOGIC_VECTOR'( and_963_nl & (NOT mux_1759_nl) & and_dcpl_837 & and_dcpl_739
      & and_965_nl));
  not_4462_nl <= NOT and_dcpl_619;
  and_966_nl <= and_dcpl_732 AND and_dcpl_826;
  nor_500_nl <= NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd OR (NOT
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1) OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("10")));
  mux_1770_nl <= MUX_s_1_2_2(mux_1555_cse, mux_1553_cse, nor_500_nl);
  mux_1772_nl <= MUX_s_1_2_2(mux_1557_cse, mux_1770_nl, fsm_output(0));
  mux_1774_nl <= MUX_s_1_2_2(mux_1559_cse, mux_1772_nl, and_1773_cse);
  mux_1775_nl <= MUX_s_1_2_2(mux_1774_nl, mux_1546_cse, fsm_output(7));
  and_968_nl <= and_dcpl_743 AND and_dcpl_740 AND and_dcpl_825;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_46_nl <= MUX1HOT_v_16_5_2(z_out_1, attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0,
      (rms_norm_16_div_cmp_z_oreg(15 DOWNTO 0)), output_0_6_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      STD_LOGIC_VECTOR'( and_966_nl & (NOT mux_1775_nl) & and_dcpl_827 & and_dcpl_739
      & and_968_nl));
  not_4461_nl <= NOT and_dcpl_619;
  and_969_nl <= and_dcpl_732 AND and_dcpl_820;
  or_2492_nl <= CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd) OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  mux_1786_nl <= MUX_s_1_2_2(mux_1553_cse, mux_1555_cse, or_2492_nl);
  mux_1788_nl <= MUX_s_1_2_2(mux_1557_cse, mux_1786_nl, fsm_output(0));
  mux_1790_nl <= MUX_s_1_2_2(mux_1559_cse, mux_1788_nl, and_1773_cse);
  mux_1791_nl <= MUX_s_1_2_2(mux_1790_nl, mux_1546_cse, fsm_output(7));
  and_971_nl <= and_dcpl_743 AND and_dcpl_551 AND and_dcpl_818;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_48_nl <= MUX1HOT_v_16_5_2(z_out_1, attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0,
      (rms_norm_16_div_cmp_z_oreg(15 DOWNTO 0)), output_0_8_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      STD_LOGIC_VECTOR'( and_969_nl & (NOT mux_1791_nl) & and_dcpl_821 & and_dcpl_739
      & and_971_nl));
  not_4460_nl <= NOT and_dcpl_619;
  and_972_nl <= and_dcpl_732 AND and_dcpl_831;
  or_2497_nl <= CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd) OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  mux_1802_nl <= MUX_s_1_2_2(mux_1553_cse, mux_1555_cse, or_2497_nl);
  mux_1804_nl <= MUX_s_1_2_2(mux_1557_cse, mux_1802_nl, fsm_output(0));
  mux_1806_nl <= MUX_s_1_2_2(mux_1559_cse, mux_1804_nl, and_1773_cse);
  mux_1807_nl <= MUX_s_1_2_2(mux_1806_nl, mux_1546_cse, fsm_output(7));
  and_974_nl <= and_dcpl_743 AND and_dcpl_551 AND and_dcpl_830;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_50_nl <= MUX1HOT_v_16_5_2(z_out_1, attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0,
      (rms_norm_16_div_cmp_z_oreg(15 DOWNTO 0)), output_0_9_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      STD_LOGIC_VECTOR'( and_972_nl & (NOT mux_1807_nl) & and_dcpl_832 & and_dcpl_739
      & and_974_nl));
  not_4459_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_68_nl <= MUX1HOT_v_8_6_2((z_out_1(15 DOWNTO
      8)), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0(15 DOWNTO 8)),
      (rms_norm_16_div_cmp_z_oreg(15 DOWNTO 8)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8,
      (output_0_2_lpi_3_15_0(15 DOWNTO 8)), (drf_output_sdt_3_sva_15_0_mx0w3(15 DOWNTO
      8)), STD_LOGIC_VECTOR'( and_1034_itm & (NOT mux_1966_itm) & and_dcpl_989 &
      and_dcpl_374 & and_dcpl_739 & and_1037_itm));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_118_nl <= MUX1HOT_v_8_6_2((z_out_1(7 DOWNTO
      0)), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0(7 DOWNTO 0)),
      (rms_norm_16_div_cmp_z_oreg(7 DOWNTO 0)), STD_LOGIC_VECTOR'( APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7
      & APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6
      & APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5
      & APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4
      & APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3
      & APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2
      & APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1
      & APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0),
      (output_0_2_lpi_3_15_0(7 DOWNTO 0)), (drf_output_sdt_3_sva_15_0_mx0w3(7 DOWNTO
      0)), STD_LOGIC_VECTOR'( and_1034_itm & (NOT mux_1966_itm) & and_dcpl_989 &
      and_dcpl_374 & and_dcpl_739 & and_1037_itm));
  not_4443_nl <= NOT and_dcpl_619;
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_39_nl <= MUX_v_24_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd
      & (reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(38 DOWNTO 16))), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(39
      DOWNTO 16)), apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_39_16, apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16,
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3(39 DOWNTO 16)), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm(39
      DOWNTO 16)), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_39_16, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_39_16,
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3(39 DOWNTO 16)), (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm(39
      DOWNTO 16)), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_39_16, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16,
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3(39 DOWNTO 16)), (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm(39
      DOWNTO 16)), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_39_16, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  attention_2_1_16_16_4_4_v_proj_re_mux1h_58_nl <= MUX1HOT_v_24_7_2(attention_2_1_16_16_4_4_v_proj_re_0_12_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_39_16,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16_mx0w1, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16_mx0w1,
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16, APPLY_ROTARY_POS_EMB_LOOP_6_mux_39_nl,
      STD_LOGIC_VECTOR'( and_dcpl_726 & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240
      & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
  not_4582_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_59_nl <= MUX1HOT_v_24_6_2(attention_2_1_16_16_4_4_v_proj_re_0_14_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16_mx0w1, apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16_mx0w1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16, STD_LOGIC_VECTOR'(
      and_dcpl_726 & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847));
  not_4583_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_60_nl <= MUX1HOT_v_24_6_2(attention_2_1_16_16_4_4_v_proj_re_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16_mx0w1, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16_mx0w1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16, STD_LOGIC_VECTOR'(
      and_dcpl_726 & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847));
  not_4584_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_61_nl <= MUX1HOT_v_24_6_2(attention_2_1_16_16_4_4_v_proj_re_0_5_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_39_16, attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16_mx0w5,
      attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_39_16, STD_LOGIC_VECTOR'( and_dcpl_726
      & and_dcpl_983 & and_dcpl_240 & and_dcpl_626 & and_dcpl_207 & and_dcpl_213));
  not_4585_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_62_nl <= MUX1HOT_v_24_6_2(attention_2_1_16_16_4_4_v_proj_re_0_6_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16_mx0w1, STD_LOGIC_VECTOR'(
      and_dcpl_726 & attention_2_1_16_16_4_4_k_proj_re_or_cse & and_dcpl_983 & and_dcpl_240
      & attention_2_1_16_16_4_4_k_proj_re_or_17_cse & and_dcpl_207));
  not_4586_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_63_nl <= MUX1HOT_v_24_6_2(attention_2_1_16_16_4_4_v_proj_re_0_8_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16, STD_LOGIC_VECTOR'( and_dcpl_726
      & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847));
  not_4587_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_64_nl <= MUX1HOT_v_24_6_2(attention_2_1_16_16_4_4_v_proj_re_0_9_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16, STD_LOGIC_VECTOR'( and_dcpl_726
      & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847));
  not_4588_nl <= NOT and_dcpl_619;
  APPLY_ROTARY_POS_EMB_LOOP_3_APPLY_ROTARY_POS_EMB_LOOP_3_nor_nl <= NOT(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_or_2_nl <= and_dcpl_1151
      OR compute_sqrt_for_i_and_2_cse;
  QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_1_nl <= MUX1HOT_s_1_6_2((LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_2(0)),
      APPLY_ROTARY_POS_EMB_LOOP_3_APPLY_ROTARY_POS_EMB_LOOP_3_nor_nl, LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0,
      GEMM_3D_FLOAT_LOOP_3_and_tmp_4_sva_mx0w2, GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_0_sva_mx0w3,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1), STD_LOGIC_VECTOR'(
      and_dcpl_725 & RMS_NORM_LOOP_2_2_i_and_9_cse & QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_or_2_nl
      & and_dcpl_1152 & and_dcpl_222 & and_dcpl_557));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_95_nl <= MUX_v_2_2_2((reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1(12
      DOWNTO 11)), STD_LOGIC_VECTOR'( "10"), and_dcpl_1363);
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_96_nl <= MUX_s_1_2_2((reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1(10)),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1, and_dcpl_1363);
  APPLY_ROTARY_POS_EMB_LOOP_6_APPLY_ROTARY_POS_EMB_LOOP_6_or_7_nl <= (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1(9))
      OR and_dcpl_1363;
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_97_nl <= MUX_s_1_2_2((reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1(8)),
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2,
      and_dcpl_1363);
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_98_nl <= MUX_v_8_2_2((reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1(7
      DOWNTO 0)), reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3,
      and_dcpl_1363);
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_99_nl <= MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_39_16,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(39 DOWNTO 16)), and_dcpl_1363);
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_100_nl <= MUX_v_8_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(15 DOWNTO 8)), and_dcpl_1363);
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_101_nl <= MUX_v_8_2_2(STD_LOGIC_VECTOR'( APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6 & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4 & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2 & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(7
      DOWNTO 0)), and_dcpl_1363);
  attention_2_1_16_16_4_4_v_proj_re_mux_nl <= MUX_v_24_2_2(output_0_7_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_63_cse);
  not_4589_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_44_nl <= MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_63_cse);
  not_4590_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_v_proj_re_mux_36_nl <= MUX_v_24_2_2(output_0_8_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_65_cse);
  not_4591_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_45_nl <= MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_65_cse);
  not_4592_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_v_proj_re_mux_37_nl <= MUX_v_24_2_2(output_0_6_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_67_cse);
  not_4593_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_46_nl <= MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_67_cse);
  not_4594_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_v_proj_re_mux_38_nl <= MUX_v_24_2_2(output_0_9_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_69_cse);
  not_4595_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_47_nl <= MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_69_cse);
  not_4596_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_v_proj_re_mux_39_nl <= MUX_v_24_2_2(output_0_5_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_71_cse);
  not_4597_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_48_nl <= MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_71_cse);
  not_4598_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_v_proj_re_mux_40_nl <= MUX_v_24_2_2(output_0_10_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_73_cse);
  not_4599_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_49_nl <= MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_73_cse);
  not_4600_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_v_proj_re_mux_41_nl <= MUX_v_24_2_2(output_0_4_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_75_cse);
  not_4601_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_50_nl <= MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_75_cse);
  not_4602_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_v_proj_re_mux_42_nl <= MUX_v_24_2_2(output_0_11_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_77_cse);
  not_4603_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_51_nl <= MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_77_cse);
  not_4604_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_v_proj_re_mux_43_nl <= MUX_v_24_2_2(output_0_3_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_79_cse);
  not_4605_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_52_nl <= MUX_v_16_2_2(apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_79_cse);
  not_4606_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_v_proj_re_mux_44_nl <= MUX_v_24_2_2(output_0_12_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_81_cse);
  not_4607_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_53_nl <= MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_81_cse);
  not_4608_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_v_proj_re_mux_45_nl <= MUX_v_24_2_2(output_0_2_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_83_cse);
  not_4609_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_54_nl <= MUX_v_16_2_2(apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_83_cse);
  not_4610_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_v_proj_re_mux_46_nl <= MUX_v_24_2_2(output_0_13_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_85_cse);
  not_4611_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_55_nl <= MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_85_cse);
  not_4612_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_v_proj_re_mux_47_nl <= MUX_v_24_2_2(output_0_1_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  not_4613_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_56_nl <= MUX_v_8_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 8)), attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  not_5055_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_60_nl <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(7)),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  attention_2_1_16_16_4_4_k_proj_re_mux_61_nl <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(6)),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  attention_2_1_16_16_4_4_k_proj_re_mux_62_nl <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(5)),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  attention_2_1_16_16_4_4_k_proj_re_mux_63_nl <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(4)),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  attention_2_1_16_16_4_4_k_proj_re_mux_64_nl <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(3)),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  attention_2_1_16_16_4_4_k_proj_re_mux_65_nl <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(2)),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  attention_2_1_16_16_4_4_k_proj_re_mux_66_nl <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(1)),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  attention_2_1_16_16_4_4_k_proj_re_mux_67_nl <= MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(0)),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  attention_2_1_16_16_4_4_v_proj_re_mux_48_nl <= MUX_v_24_2_2(output_0_14_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_89_cse);
  not_4615_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_57_nl <= MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_89_cse);
  not_4616_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_v_proj_re_mux_49_nl <= MUX_v_24_2_2(output_0_0_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_91_cse);
  not_4617_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_58_nl <= MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_91_cse);
  not_4618_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_v_proj_re_mux_50_nl <= MUX_v_24_2_2(output_0_15_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(39
      DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_re_and_93_cse);
  not_4619_nl <= NOT and_dcpl_1154;
  attention_2_1_16_16_4_4_k_proj_re_mux_59_nl <= MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_re_and_93_cse);
  not_4620_nl <= NOT and_dcpl_1154;
  GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_4_nl <= NOT(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva_mx0w0
      AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  GEMM_3D_FLOAT_LOOP_3_1_and_32_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_4_nl);
  GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_6_nl <= NOT(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva_mx0w0
      AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  GEMM_3D_FLOAT_LOOP_3_1_and_34_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_6_nl);
  GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_2_nl <= NOT(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva_mx0w0
      AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  GEMM_3D_FLOAT_LOOP_3_1_and_30_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_2_nl);
  GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_12_nl <= NOT(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_1_sva_mx0w3
      AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  GEMM_3D_FLOAT_LOOP_3_1_and_40_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_12_nl);
  GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_10_nl <= NOT(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva_mx0w3
      AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  GEMM_3D_FLOAT_LOOP_3_1_and_38_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_10_nl);
  GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_14_nl <= NOT(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_0_sva_mx0w3
      AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  GEMM_3D_FLOAT_LOOP_3_1_and_42_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_14_nl);
  mux_789_nl <= MUX_s_1_2_2((NOT or_tmp_704), and_1651_cse, fsm_output(7));
  and_259_nl <= mux_789_nl AND and_dcpl_226 AND nor_1026_cse AND and_dcpl;
  and_267_nl <= and_dcpl_185 AND nor_777_cse AND (NOT (fsm_output(5))) AND and_dcpl_231
      AND (fsm_output(7)) AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd) AND
      LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0;
  or_1734_nl <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd OR (NOT(LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11"))));
  mux_793_nl <= MUX_s_1_2_2(mux_792_cse, or_1734_nl, fsm_output(3));
  mux_794_nl <= MUX_s_1_2_2(mux_793_nl, or_tmp_708, fsm_output(2));
  nand_307_nl <= NOT((fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(7)));
  mux_791_nl <= MUX_s_1_2_2(or_tmp_708, nand_307_nl, fsm_output(2));
  mux_795_nl <= MUX_s_1_2_2(mux_794_nl, mux_791_nl, or_1732_cse);
  nand_308_nl <= NOT(((fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(6))) AND
      (fsm_output(7)));
  nand_309_nl <= NOT(((NOT (fsm_output(1))) OR (fsm_output(2)) OR (fsm_output(3))
      OR (fsm_output(6))) AND (fsm_output(7)));
  mux_790_nl <= MUX_s_1_2_2(nand_308_nl, nand_309_nl, fsm_output(0));
  mux_796_nl <= MUX_s_1_2_2(mux_795_nl, mux_790_nl, fsm_output(4));
  mux_797_nl <= MUX_s_1_2_2(mux_796_nl, (NOT (fsm_output(7))), fsm_output(5));
  nor_980_nl <= NOT((fsm_output(1)) OR (fsm_output(8)));
  nor_981_nl <= NOT((fsm_output(1)) OR (fsm_output(0)) OR (fsm_output(8)));
  or_1854_nl <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd OR (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1))
      OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 OR (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0));
  mux_897_nl <= MUX_s_1_2_2(nor_980_nl, nor_981_nl, or_1854_nl);
  mux_898_nl <= MUX_s_1_2_2(mux_897_nl, (fsm_output(8)), fsm_output(5));
  mux_899_nl <= MUX_s_1_2_2(mux_898_nl, nor_tmp_307, fsm_output(3));
  mux_896_nl <= MUX_s_1_2_2(nor_tmp_307, (fsm_output(5)), fsm_output(3));
  mux_900_nl <= MUX_s_1_2_2(mux_899_nl, mux_896_nl, fsm_output(4));
  or_1857_nl <= (fsm_output(6)) OR mux_900_nl;
  and_380_nl <= (fsm_output(5)) AND (and_1474_cse OR (fsm_output(8)));
  mux_894_nl <= MUX_s_1_2_2(and_380_nl, or_1851_cse, fsm_output(3));
  mux_895_nl <= MUX_s_1_2_2(nor_tmp_307, mux_894_nl, fsm_output(4));
  or_1853_nl <= (fsm_output(6)) OR mux_895_nl;
  mux_901_nl <= MUX_s_1_2_2(or_1857_nl, or_1853_nl, fsm_output(2));
  nand_316_nl <= NOT((fsm_output(3)) AND (fsm_output(5)) AND (fsm_output(1)) AND
      (NOT (fsm_output(8))));
  or_1849_nl <= (fsm_output(3)) OR (fsm_output(5)) OR (NOT (fsm_output(1))) OR (NOT
      (fsm_output(0))) OR (fsm_output(8));
  mux_891_nl <= MUX_s_1_2_2(nand_316_nl, or_1849_nl, fsm_output(4));
  mux_888_nl <= MUX_s_1_2_2(or_1848_cse, (fsm_output(8)), fsm_output(5));
  or_1847_nl <= nor_305_cse OR (fsm_output(8));
  mux_889_nl <= MUX_s_1_2_2(mux_888_nl, or_1847_nl, fsm_output(3));
  mux_890_nl <= MUX_s_1_2_2(mux_889_nl, (fsm_output(8)), fsm_output(4));
  mux_892_nl <= MUX_s_1_2_2(mux_891_nl, mux_890_nl, fsm_output(6));
  or_1846_nl <= (NOT (fsm_output(4))) OR (fsm_output(3)) OR (fsm_output(5)) OR (fsm_output(1))
      OR (fsm_output(0)) OR (fsm_output(8));
  or_1845_nl <= (NOT(CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)/=STD_LOGIC_VECTOR'("00")) OR reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 OR
      (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0)) OR (NOT (fsm_output(4))) OR (fsm_output(3))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(0)))))
      OR (fsm_output(8));
  mux_887_nl <= MUX_s_1_2_2(or_1846_nl, or_1845_nl, fsm_output(6));
  mux_893_nl <= MUX_s_1_2_2(mux_892_nl, mux_887_nl, fsm_output(2));
  mux_902_nl <= MUX_s_1_2_2(mux_901_nl, mux_893_nl, fsm_output(7));
  GEMM_3D_FLOAT_LOOP_4_1_mux_17_nl <= MUX_s_1_16_2((apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2(39)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2(39)), (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2(39)),
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2(39)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2(39)), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2(39)),
      (attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3(39)), (attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3(39)),
      (attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3(39)), (attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3(39)),
      (attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3(39)), (attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3(39)),
      (attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3(39)), (attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3(39)),
      (attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3(39)), STD_LOGIC_VECTOR'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1));
  rms_norm_16_variance_mux1h_nl <= MUX1HOT_s_1_9_2((acc_3_cse_40_1(39)), (compute_sqrt_for_acc_1_itm_40_1_1(39)),
      attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_39, (APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1(39)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux1h_5_itm(39)), (softmax_1_4_3_sum_sva_2(39)), (SOFTMAX_LOOP_5_mux_12_psp_mx0w0(39)),
      GEMM_3D_FLOAT_LOOP_4_1_mux_17_nl, (compute_sqrt_1_for_acc_1_itm_40_1_1(39)),
      STD_LOGIC_VECTOR'( rms_norm_16_variance_or_1_cse & and_dcpl_290 & and_404_itm
      & and_dcpl_374 & and_dcpl_313 & and_dcpl_377 & and_dcpl_294 & and_dcpl_316
      & and_dcpl_292));
  GEMM_3D_FLOAT_LOOP_4_1_mux_24_nl <= MUX_v_39_16_2((apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2(38
      DOWNTO 0)), (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2(38 DOWNTO 0)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2(38 DOWNTO 0)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1,
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2(38 DOWNTO 0)), (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2(38
      DOWNTO 0)), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2(38 DOWNTO 0)),
      (attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3(38 DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3(38
      DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3(38 DOWNTO 0)),
      (attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3(38 DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3(38
      DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3(38 DOWNTO 0)),
      (attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3(38 DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3(38
      DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3(38 DOWNTO 0)),
      STD_LOGIC_VECTOR'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1));
  rms_norm_16_variance_mux1h_1_nl <= MUX1HOT_v_39_10_2((acc_3_cse_40_1(38 DOWNTO
      0)), (compute_sqrt_for_acc_1_itm_40_1_1(38 DOWNTO 0)), (attention_abs_1_qr_sva_1(38
      DOWNTO 0)), attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_38_0,
      (APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1(38 DOWNTO 0)), (GEMM_3D_FLOAT_LOOP_4_1_mux1h_5_itm(38
      DOWNTO 0)), (softmax_1_4_3_sum_sva_2(38 DOWNTO 0)), (SOFTMAX_LOOP_5_mux_12_psp_mx0w0(38
      DOWNTO 0)), GEMM_3D_FLOAT_LOOP_4_1_mux_24_nl, (compute_sqrt_1_for_acc_1_itm_40_1_1(38
      DOWNTO 0)), STD_LOGIC_VECTOR'( rms_norm_16_variance_or_1_cse & and_dcpl_290
      & and_dcpl_363 & and_404_itm & and_dcpl_374 & and_dcpl_313 & and_dcpl_377 &
      and_dcpl_294 & and_dcpl_316 & and_dcpl_292));
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux_nl <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0(3)),
      (z_out_12(3)), LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_cse);
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_8_nl <= MUX1HOT_s_1_5_2((LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0(2)),
      (z_out_12(2)), (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_15_sdt_1(2)), (z_out_3(2)),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1, STD_LOGIC_VECTOR'(
      and_416_itm & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_cse & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_7_cse
      & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_8_cse & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_9_cse));
  and_1238_nl <= nor_1314_cse AND and_dcpl_200 AND and_dcpl_885;
  QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux_nl <= MUX_v_2_2_2(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2,
      (z_out_3(1 DOWNTO 0)), and_1238_nl);
  mux_2231_nl <= MUX_s_1_2_2((NOT nor_tmp_329), or_tmp_1221, fsm_output(3));
  mux_2230_nl <= MUX_s_1_2_2(or_tmp_992, or_tmp_861, fsm_output(3));
  mux_2232_nl <= MUX_s_1_2_2(mux_2231_nl, mux_2230_nl, fsm_output(6));
  nor_1322_nl <= NOT(mux_2232_nl OR or_1851_cse OR (NOT (fsm_output(7))));
  QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_1_nl
      <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux_nl,
      nor_1322_nl);
  nor_996_nl <= NOT(and_1474_cse OR (fsm_output(2)) OR (NOT (fsm_output(4))));
  mux_983_nl <= MUX_s_1_2_2(and_1570_cse, nor_996_nl, fsm_output(3));
  mux_982_nl <= MUX_s_1_2_2(or_270_cse, or_tmp_861, fsm_output(3));
  mux_984_nl <= MUX_s_1_2_2(mux_983_nl, (NOT mux_982_nl), fsm_output(6));
  and_426_nl <= mux_984_nl AND and_dcpl_388;
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_9_nl <= MUX1HOT_v_2_6_2((LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0(1
      DOWNTO 0)), (z_out_12(1 DOWNTO 0)), QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_1_nl,
      (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_15_sdt_1(1 DOWNTO 0)), (z_out_3(1 DOWNTO
      0)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2, STD_LOGIC_VECTOR'(
      and_416_itm & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_cse & and_426_nl & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_7_cse
      & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_8_cse & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_9_cse));
  compute_sqrt_for_i_mux1h_nl <= MUX1HOT_s_1_4_2((LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1(3)),
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp(3)), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0(3)),
      (RMS_NORM_LOOP_2_2_i_4_0_sva_1(3)), STD_LOGIC_VECTOR'( and_dcpl_242 & LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c2
      & LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c5 & and_dcpl_410));
  compute_sqrt_for_i_mux1h_1_nl <= MUX1HOT_v_2_7_2((LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1(2
      DOWNTO 1)), (LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp(2 DOWNTO 1)), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0(2
      DOWNTO 1)), (RMS_NORM_LOOP_2_2_i_4_0_sva_1(2 DOWNTO 1)), (z_out_5(2 DOWNTO
      1)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1, (z_out_11(2 DOWNTO
      1)), STD_LOGIC_VECTOR'( and_dcpl_242 & LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c2
      & LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c5 & and_dcpl_410 & compute_sqrt_for_i_and_cse
      & compute_sqrt_for_i_and_4_cse & compute_sqrt_for_i_and_5_cse));
  LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_not_2_nl <= NOT LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c3;
  compute_sqrt_for_i_nand_1_nl <= NOT(MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), compute_sqrt_for_i_mux1h_1_nl,
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_not_2_nl));
  compute_sqrt_for_i_or_nl <= compute_sqrt_for_i_and_4_cse OR compute_sqrt_for_i_and_2_cse;
  compute_sqrt_for_i_mux1h_2_nl <= MUX1HOT_s_1_8_2((LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1(0)),
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp(0)), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0(0)),
      (RMS_NORM_LOOP_2_2_i_4_0_sva_1(0)), (z_out_5(0)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2,
      (z_out_11(0)), (NOT QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1),
      STD_LOGIC_VECTOR'( and_dcpl_242 & LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c2
      & LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c5 & and_dcpl_410 & compute_sqrt_for_i_and_cse
      & compute_sqrt_for_i_or_nl & compute_sqrt_for_i_and_5_cse & and_dcpl_557));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_37_nl <= MUX_s_1_16_2(QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39,
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd, (apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_39_16(23)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16(23)), (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3(39)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm(39)), (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_39_16(23)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16(23)), (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3(39)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm(39)), (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_39_16(23)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16(23)), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3(39)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm(39)), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_39_16(23)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16(23)), STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_69_nl <= MUX_v_23_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(38
      DOWNTO 16)), (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1(38 DOWNTO
      16)), (apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_39_16(22 DOWNTO 0)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16(22 DOWNTO 0)), (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3(38
      DOWNTO 16)), (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm(38 DOWNTO
      16)), (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_39_16(22 DOWNTO 0)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16(22 DOWNTO 0)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3(38 DOWNTO 16)), (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm(38
      DOWNTO 16)), (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_39_16(22 DOWNTO
      0)), (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16(22 DOWNTO
      0)), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3(38 DOWNTO 16)), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm(38
      DOWNTO 16)), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_39_16(22 DOWNTO
      0)), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16(22 DOWNTO
      0)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd &
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  nand_373_nl <= NOT((reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 OR (NOT reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1)
      OR reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 OR reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd)
      AND (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(1)) AND (fsm_output(0))
      AND (NOT (fsm_output(6))) AND (fsm_output(7)));
  nor_576_nl <= NOT((NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      OR (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1))) OR CONV_SL_1_1(fsm_output(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")));
  mux_2079_nl <= MUX_s_1_2_2(or_1983_cse, mux_806_cse, nor_576_nl);
  mux_2080_nl <= MUX_s_1_2_2(nand_373_nl, mux_2079_nl, fsm_output(4));
  or_2775_nl <= (fsm_output(1)) OR (fsm_output(0)) OR (NOT (fsm_output(6))) OR (fsm_output(7));
  mux_2077_nl <= MUX_s_1_2_2(or_1983_cse, or_2775_nl, and_1773_cse);
  or_2777_nl <= (fsm_output(4)) OR mux_2077_nl;
  mux_2081_nl <= MUX_s_1_2_2(mux_2080_nl, or_2777_nl, fsm_output(5));
  nor_1225_nl <= NOT(mux_2081_nl OR (fsm_output(8)));
  and_1110_nl <= and_dcpl_1061 AND and_dcpl_45 AND (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd)
      AND (NOT(reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 OR reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0))
      AND reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  and_1115_nl <= and_dcpl_205 AND and_dcpl_421 AND and_dcpl_319 AND (NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd)) AND reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  INIT_2D_MEM_LOOP_2_1_mux1h_nl <= MUX1HOT_v_24_9_2(attention_2_1_16_16_4_4_v_proj_re_0_10_sva_1_39_16,
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_conc_1_mut_71_48_mx0w0, for_for_strm_in_tmp_sva_25_2,
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_39_16,
      RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_39_16, APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1,
      (APPLY_ROTARY_POS_EMB_LOOP_6_mux_37_nl & APPLY_ROTARY_POS_EMB_LOOP_6_mux_69_nl),
      STD_LOGIC_VECTOR'( and_dcpl_726 & and_dcpl_257 & nor_1225_nl & and_dcpl_1011
      & and_dcpl_983 & and_1110_nl & and_dcpl_847 & and_1115_nl & and_dcpl_583));
  mux_2074_nl <= MUX_s_1_2_2((NOT or_tmp_728), or_tmp_767, fsm_output(5));
  mux_2075_nl <= MUX_s_1_2_2(mux_tmp_91, mux_2074_nl, fsm_output(3));
  nand_96_nl <= NOT((fsm_output(6)) AND (NOT mux_2075_nl));
  mux_2076_nl <= MUX_s_1_2_2(nand_96_nl, or_tmp_913, fsm_output(7));
  nor_1323_nl <= NOT(mux_2076_nl OR (fsm_output(8)));
  INIT_2D_MEM_LOOP_2_1_and_nl <= MUX_v_24_2_2(STD_LOGIC_VECTOR'("000000000000000000000000"),
      INIT_2D_MEM_LOOP_2_1_mux1h_nl, nor_1323_nl);
  GEMM_3D_FLOAT_LOOP_4_mux_17_nl <= MUX_v_40_16_2(attention_2_1_16_16_4_4_q_embed_0_0_0_sva_1,
      attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1, attention_2_1_16_16_4_4_q_embed_0_0_2_sva_1,
      attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1, attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1,
      attention_2_1_16_16_4_4_q_embed_1_0_1_sva_1, attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1,
      attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1, attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1,
      attention_2_1_16_16_4_4_q_embed_2_0_1_sva_1, attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1,
      attention_2_1_16_16_4_4_q_embed_2_0_3_sva_1, attention_2_1_16_16_4_4_q_embed_3_0_0_sva_1,
      attention_2_1_16_16_4_4_q_embed_3_0_1_sva_1, attention_2_1_16_16_4_4_q_embed_3_0_2_sva_1,
      attention_2_1_16_16_4_4_q_embed_3_0_3_sva_1, STD_LOGIC_VECTOR'( reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1));
  SOFTMAX_LOOP_4_x_mux_nl <= MUX_v_40_12_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9,
      attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9, attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9,
      attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9, attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8,
      attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8, attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8,
      attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8, attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8,
      attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8, attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8,
      attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1));
  SOFTMAX_LOOP_4_x_acc_2_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(SOFTMAX_LOOP_4_x_mux_nl)
      + SIGNED((NOT QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39) & (NOT
      QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0)) + SIGNED'( "0000000000000000000000000000000000000001"),
      40));
  GEMM_3D_FLOAT_LOOP_4_1_mux_18_nl <= MUX_v_40_12_2(attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1, reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  mux_1059_nl <= MUX_s_1_2_2(or_tmp_930, mux_tmp_1044, fsm_output(1));
  mux_1058_nl <= MUX_s_1_2_2(or_tmp_930, or_tmp_931, fsm_output(1));
  mux_1060_nl <= MUX_s_1_2_2(mux_1059_nl, mux_1058_nl, fsm_output(0));
  mux_1057_nl <= MUX_s_1_2_2(mux_tmp_1051, or_tmp_930, fsm_output(1));
  mux_1061_nl <= MUX_s_1_2_2(mux_1060_nl, mux_1057_nl, fsm_output(3));
  mux_1054_nl <= MUX_s_1_2_2(or_tmp_931, mux_tmp_1052, fsm_output(1));
  mux_1053_nl <= MUX_s_1_2_2(mux_tmp_1052, mux_tmp_1051, fsm_output(1));
  mux_1055_nl <= MUX_s_1_2_2(mux_1054_nl, mux_1053_nl, fsm_output(0));
  or_1996_nl <= (fsm_output(1)) OR (fsm_output(4)) OR (NOT (fsm_output(7)));
  mux_1050_nl <= MUX_s_1_2_2(or_tmp_930, or_1996_nl, fsm_output(0));
  mux_1056_nl <= MUX_s_1_2_2(mux_1055_nl, mux_1050_nl, fsm_output(3));
  mux_1062_nl <= MUX_s_1_2_2(mux_1061_nl, mux_1056_nl, fsm_output(2));
  or_1994_nl <= nor_646_cse OR (fsm_output(7));
  mux_1047_nl <= MUX_s_1_2_2((NOT mux_tmp_1044), (fsm_output(7)), or_1732_cse);
  mux_1048_nl <= MUX_s_1_2_2(or_1994_nl, mux_1047_nl, fsm_output(3));
  mux_1042_nl <= MUX_s_1_2_2((fsm_output(7)), (NOT (fsm_output(7))), fsm_output(4));
  mux_1043_nl <= MUX_s_1_2_2(mux_1042_nl, or_tmp_922, fsm_output(5));
  mux_1045_nl <= MUX_s_1_2_2(mux_tmp_1044, mux_1043_nl, nor_366_cse);
  mux_1046_nl <= MUX_s_1_2_2((NOT mux_1045_nl), (fsm_output(7)), fsm_output(3));
  mux_1049_nl <= MUX_s_1_2_2(mux_1048_nl, mux_1046_nl, fsm_output(2));
  mux_1063_nl <= MUX_s_1_2_2(mux_1062_nl, mux_1049_nl, fsm_output(6));
  RMS_NORM_LOOP_2_mux_22_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1(39)),
      (input_0_1_sva_1(39)), input_0_2_sva_1_39, (input_0_3_sva_1(39)), (input_0_4_sva_1(39)),
      (input_0_5_sva_1(39)), (input_0_6_sva_1(39)), (input_0_7_sva_1(39)), (input_0_8_sva_1(39)),
      (input_0_9_sva_1(39)), (input_0_10_sva_1(39)), (input_0_11_sva_1(39)), (input_0_12_sva_1(39)),
      input_0_13_sva_1_39, (input_0_14_sva_1(39)), (attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3(39)),
      reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  QUANTIZE_ACTIVATION_LOOP_3_quantized_value_mux_nl <= MUX_s_1_16_2((input_0_0_sva_2(39)),
      (input_0_1_sva_2(39)), input_0_2_sva_2_39, (input_0_3_sva_2(39)), (input_0_4_sva_2(39)),
      (input_0_5_sva_2(39)), (input_0_6_sva_2(39)), (input_0_7_sva_2(39)), (input_0_8_sva_2(39)),
      (input_0_9_sva_2(39)), (input_0_10_sva_2(39)), (input_0_11_sva_2(39)), (input_0_12_sva_2(39)),
      input_0_13_sva_2_39, (input_0_14_sva_2(39)), (input_0_15_sva_1(39)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  RMS_NORM_LOOP_2_mux_24_nl <= MUX_v_39_16_2((attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1(38
      DOWNTO 0)), (input_0_1_sva_1(38 DOWNTO 0)), input_0_2_sva_1_38_0, (input_0_3_sva_1(38
      DOWNTO 0)), (input_0_4_sva_1(38 DOWNTO 0)), (input_0_5_sva_1(38 DOWNTO 0)),
      (input_0_6_sva_1(38 DOWNTO 0)), (input_0_7_sva_1(38 DOWNTO 0)), (input_0_8_sva_1(38
      DOWNTO 0)), (input_0_9_sva_1(38 DOWNTO 0)), (input_0_10_sva_1(38 DOWNTO 0)),
      (input_0_11_sva_1(38 DOWNTO 0)), (input_0_12_sva_1(38 DOWNTO 0)), input_0_13_sva_1_38_0,
      (input_0_14_sva_1(38 DOWNTO 0)), (attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3(38
      DOWNTO 0)), reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  QUANTIZE_ACTIVATION_LOOP_3_quantized_value_mux_1_nl <= MUX_v_39_16_2((input_0_0_sva_2(38
      DOWNTO 0)), (input_0_1_sva_2(38 DOWNTO 0)), input_0_2_sva_2_38_0, (input_0_3_sva_2(38
      DOWNTO 0)), (input_0_4_sva_2(38 DOWNTO 0)), (input_0_5_sva_2(38 DOWNTO 0)),
      (input_0_6_sva_2(38 DOWNTO 0)), (input_0_7_sva_2(38 DOWNTO 0)), (input_0_8_sva_2(38
      DOWNTO 0)), (input_0_9_sva_2(38 DOWNTO 0)), (input_0_10_sva_2(38 DOWNTO 0)),
      (input_0_11_sva_2(38 DOWNTO 0)), (input_0_12_sva_2(38 DOWNTO 0)), input_0_13_sva_2_38_0,
      (input_0_14_sva_2(38 DOWNTO 0)), (input_0_15_sva_1(38 DOWNTO 0)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  for_for_for_for_nand_nl <= NOT(mux_1079_itm AND (NOT(or_dcpl_1025 AND and_dcpl_204)));
  for_for_and_24_nl <= (NOT or_dcpl_1025) AND and_dcpl_204;
  for_for_mux1h_5_nl <= MUX1HOT_v_40_9_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),40)),
      input_0_12_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1, APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_q_embed_0_0_0_sva_1, attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2,
      attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx2, (ATTN_2D_LOOP_3_mux_16_itm
      & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c0 &
      attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c1 & for_for_for_for_nand_nl
      & for_for_and_24_nl & and_dcpl_216 & and_dcpl_348 & and_dcpl_351 & and_dcpl_352
      & attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c9));
  attention_2_1_16_16_4_4_attn_output_2D_not_nl <= NOT attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c7;
  for_for_mux1h_6_nl <= MUX1HOT_v_40_8_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),40)),
      input_0_7_sva_1, attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1, attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1_mx0w1,
      attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2, attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx1,
      (ATTN_2D_LOOP_3_mux_16_itm & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c0
      & attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c1 & and_dcpl_346 &
      and_dcpl_204 & and_dcpl_348 & and_dcpl_351 & and_dcpl_352 & attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c9));
  attention_2_1_16_16_4_4_attn_output_2D_not_3_nl <= NOT attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c7;
  or_2048_nl <= (NOT(CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)/=STD_LOGIC_VECTOR'("10")) OR reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 OR
      (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0))) OR CONV_SL_1_1(fsm_output(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10111")))) OR (fsm_output(8));
  mux_1095_nl <= MUX_s_1_2_2(mux_1074_cse, or_2048_nl, fsm_output(5));
  mux_1097_nl <= MUX_s_1_2_2(nand_50_cse, mux_1095_nl, fsm_output(6));
  mux_1099_nl <= MUX_s_1_2_2(or_2029_cse, mux_1097_nl, fsm_output(7));
  GEMM_3D_FLOAT_LOOP_3_1_and_36_nl <= reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd
      AND GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_8_seb;
  GEMM_3D_FLOAT_LOOP_3_1_and_52_nl <= MUX_v_39_2_2(STD_LOGIC_VECTOR'("000000000000000000000000000000000000000"),
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_8_seb);
  for_for_and_22_nl <= (NOT and_dcpl_548) AND and_dcpl_477;
  GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_nl <= NOT(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva_mx0w0
      AND (NOT reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  GEMM_3D_FLOAT_LOOP_3_1_and_28_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_nl);
  and_521_nl <= and_dcpl_342 AND and_dcpl_336 AND and_dcpl_480;
  and_523_nl <= or_dcpl_1084 AND and_dcpl_185 AND and_dcpl_422;
  GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_1_nl <= NOT(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_0_sva_mx0w3
      AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd);
  GEMM_3D_FLOAT_LOOP_3_1_and_29_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_1_nl);
  and_527_nl <= and_dcpl_342 AND and_dcpl_417 AND and_dcpl_486;
  and_529_nl <= or_dcpl_1085 AND and_dcpl_185 AND and_dcpl_422;
  GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_3_nl <= NOT(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_1_sva_mx0w3
      AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd);
  GEMM_3D_FLOAT_LOOP_3_1_and_31_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_3_nl);
  and_531_nl <= and_dcpl_342 AND and_dcpl_336 AND and_dcpl_486;
  and_533_nl <= or_dcpl_1086 AND and_dcpl_185 AND and_dcpl_422;
  GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_5_nl <= NOT(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva_mx0w3
      AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd);
  GEMM_3D_FLOAT_LOOP_3_1_and_33_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_5_nl);
  and_535_nl <= and_dcpl_342 AND and_dcpl_417 AND and_dcpl_480;
  and_537_nl <= or_dcpl_1087 AND and_dcpl_185 AND and_dcpl_422;
  GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_7_nl <= NOT(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva_mx0w3
      AND reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd);
  GEMM_3D_FLOAT_LOOP_3_1_and_35_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_7_nl);
  and_539_nl <= and_dcpl_342 AND and_dcpl_336 AND and_dcpl_471;
  and_541_nl <= or_dcpl_1088 AND and_dcpl_185 AND and_dcpl_422;
  for_for_or_4_nl <= attention_2_1_16_16_4_4_q_embed_and_24_cse OR and_dcpl_222 OR
      (nand_302_cse AND and_dcpl_187);
  for_for_and_28_nl <= (NOT nand_302_cse) AND and_dcpl_187;
  for_for_mux1h_13_nl <= MUX1HOT_v_40_8_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),40)),
      input_0_10_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_3_sva_1, APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3, acc_3_cse_40_1, (ATTN_2D_LOOP_3_mux_16_itm
      & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c0 &
      attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c1 & and_dcpl_346 & attention_2_1_16_16_4_4_q_embed_and_23_cse
      & for_for_or_4_nl & for_for_and_28_nl & and_dcpl_352 & attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c10));
  for_for_or_3_nl <= MUX_v_40_2_2(for_for_mux1h_13_nl, STD_LOGIC_VECTOR'("1111111111111111111111111111111111111111"),
      attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c8);
  or_nl <= ((NOT (z_out_5(2))) AND attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c8)
      OR attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c5;
  mux_nl <= MUX_v_40_2_2(for_for_or_3_nl, attention_2_1_16_16_4_4_attn_output_3_0_0_sva_2,
      or_nl);
  nor_nl <= NOT((GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva_mx0w0 AND and_dcpl_222 AND
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd) OR ((z_out_5(2)) AND attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c8));
  or_2087_nl <= (NOT(CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)/=STD_LOGIC_VECTOR'("11")) OR reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 OR
      (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0)) OR CONV_SL_1_1(fsm_output(4 DOWNTO
      0)/=STD_LOGIC_VECTOR'("10111")))) OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011"));
  mux_1133_nl <= MUX_s_1_2_2(mux_1132_cse, or_2087_nl, fsm_output(5));
  or_3215_nl <= (NOT mux_1147_itm) OR (and_dcpl_222 AND (NOT or_3212_tmp)) OR attention_2_1_16_16_4_4_attn_output_and_14_cse
      OR attention_2_1_16_16_4_4_q_embed_and_26_cse;
  mux1h_nl <= MUX1HOT_v_40_9_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),40)),
      input_0_4_sva_1, attention_2_1_16_16_4_4_k_embed_3_0_0_sva_1, attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1, attention_2_1_16_16_4_4_attn_output_3_0_1_sva_2,
      acc_3_cse_40_1, (ATTN_2D_LOOP_3_mux_16_itm & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c0 &
      attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c1 & and_dcpl_346 & or_3215_nl
      & attention_2_1_16_16_4_4_q_embed_and_25_cse & and_dcpl_524 & attention_2_1_16_16_4_4_attn_output_and_13_cse
      & and_dcpl_352 & attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c10));
  not_4622_nl <= NOT or_3212_tmp;
  or_3216_nl <= (NOT mux_1177_itm) OR (and_dcpl_222 AND (NOT or_3213_tmp)) OR attention_2_1_16_16_4_4_attn_output_and_16_cse
      OR attention_2_1_16_16_4_4_q_embed_and_28_cse;
  mux1h_1_nl <= MUX1HOT_v_40_9_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),40)),
      input_0_11_sva_1, attention_2_1_16_16_4_4_k_embed_3_0_1_sva_1, attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1, attention_2_1_16_16_4_4_attn_output_3_0_2_sva_2,
      acc_3_cse_40_1, (ATTN_2D_LOOP_3_mux_16_itm & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c0 &
      attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c1 & and_dcpl_346 & or_3216_nl
      & attention_2_1_16_16_4_4_q_embed_and_27_cse & and_dcpl_524 & attention_2_1_16_16_4_4_attn_output_and_15_cse
      & and_dcpl_352 & attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c10));
  not_4624_nl <= NOT or_3213_tmp;
  or_3217_nl <= (NOT mux_1197_itm) OR (and_dcpl_222 AND (NOT or_3214_tmp)) OR attention_2_1_16_16_4_4_attn_output_and_18_cse
      OR attention_2_1_16_16_4_4_q_embed_and_30_cse;
  mux1h_2_nl <= MUX1HOT_v_40_11_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(strm_in_rsci_idat_mxwt),40)),
      input_0_3_sva_1, STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(for_for_strm_in_tmp_sva_31_26
      & for_for_strm_in_tmp_sva_25_2),40)), attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3,
      input_0_15_sva_1, attention_2_1_16_16_4_4_k_embed_3_0_2_sva_1, APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_3_0_3_sva_2, acc_3_cse_40_1, (ATTN_2D_LOOP_3_mux_16_itm
      & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c0 &
      attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c1 & and_dcpl_242 & or_3217_nl
      & and_dcpl_344 & and_dcpl_346 & attention_2_1_16_16_4_4_q_embed_and_29_cse
      & and_dcpl_524 & attention_2_1_16_16_4_4_attn_output_and_17_cse & and_dcpl_352
      & attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c12));
  not_4626_nl <= NOT or_3214_tmp;
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_7_nl <= MUX1HOT_s_1_5_2((z_out_12(4)), (compute_sqrt_for_acc_1_itm_40_1_1(39)),
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp(4)), (compute_sqrt_1_for_acc_1_itm_40_1_1(39)),
      (RMS_NORM_LOOP_2_2_acc_1_tmp(4)), STD_LOGIC_VECTOR'( and_581_ssc & and_dcpl_290
      & and_dcpl_439 & and_dcpl_292 & and_dcpl_306));
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_10_nl <= MUX1HOT_v_4_6_2((z_out_12(3 DOWNTO
      0)), (compute_sqrt_for_acc_1_itm_40_1_1(38 DOWNTO 35)), (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2),
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp(3 DOWNTO 0)), (compute_sqrt_1_for_acc_1_itm_40_1_1(38
      DOWNTO 35)), (RMS_NORM_LOOP_2_2_acc_1_tmp(3 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_581_ssc & and_dcpl_290 & and_dcpl_477 & and_dcpl_439 & and_dcpl_292 & and_dcpl_306));
  LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_4_nl <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"),
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_10_nl, LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_nand_seb);
  attention_2_1_16_16_4_4_q_proj_attention_2_1_16_16_4_4_q_proj_mux_12_nl <= MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_15,
      (z_out(15)), and_1191_rgt);
  operator_40_24_true_AC_TRN_AC_WRAP_1_and_2_nl <= (NOT and_dcpl_739) AND (NOT mux_1309_cse)
      AND (fsm_output(2)) AND and_dcpl_577 AND and_dcpl_576;
  RMS_NORM_LOOP_2_2_i_mux1h_3_nl <= MUX1HOT_v_3_3_2((RMS_NORM_LOOP_2_2_i_4_0_sva_1(3
      DOWNTO 1)), (LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1(3 DOWNTO 1)), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0(3
      DOWNTO 1)), STD_LOGIC_VECTOR'( and_dcpl_477 & and_dcpl_410 & and_dcpl_255));
  RMS_NORM_LOOP_2_2_i_not_2_nl <= NOT RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c1;
  APPLY_ROTARY_POS_EMB_LOOP_3_and_10_nl <= reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      AND (NOT reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  RMS_NORM_LOOP_2_2_i_mux1h_6_nl <= MUX1HOT_s_1_7_2((RMS_NORM_LOOP_2_2_i_4_0_sva_1(0)),
      (LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1(0)), APPLY_ROTARY_POS_EMB_LOOP_3_and_10_nl,
      GEMM_3D_FLOAT_LOOP_3_and_tmp_5_sva_mx0w2, GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_1_sva_mx0w3,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0(0)),
      STD_LOGIC_VECTOR'( and_dcpl_477 & and_dcpl_410 & RMS_NORM_LOOP_2_2_i_and_9_cse
      & and_dcpl_1152 & and_dcpl_222 & and_dcpl_557 & and_dcpl_255));
  or_2335_nl <= and_1638_cse OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_1433_nl <= MUX_s_1_2_2(or_2335_nl, or_1983_cse, fsm_output(5));
  mux_1428_nl <= MUX_s_1_2_2(or_1983_cse, (NOT (fsm_output(6))), fsm_output(0));
  nor_1105_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  mux_1429_nl <= MUX_s_1_2_2(mux_1428_nl, nor_1105_nl, fsm_output(1));
  mux_1430_nl <= MUX_s_1_2_2(or_1983_cse, mux_1429_nl, fsm_output(2));
  or_2331_nl <= (NOT(nor_1106_cse OR (fsm_output(6)))) OR (fsm_output(7));
  mux_1431_nl <= MUX_s_1_2_2(mux_1430_nl, or_2331_nl, fsm_output(3));
  mux_1432_nl <= MUX_s_1_2_2(or_1983_cse, mux_1431_nl, fsm_output(5));
  mux_1434_nl <= MUX_s_1_2_2(mux_1433_nl, mux_1432_nl, fsm_output(4));
  QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_nl <= MUX1HOT_s_1_3_2(reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0,
      (z_out_3(1)), (z_out_3(1)), STD_LOGIC_VECTOR'( QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_or_cse
      & and_dcpl_726 & and_937_ssc));
  QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_3_nl <= QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_nl
      AND nor_1324_seb;
  RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_and_nl <= (LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp(4))
      AND RMS_NORM_LOOP_2_2_unequal_tmp_mx0w0;
  QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_3_nl <= MUX1HOT_s_1_3_2(reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1,
      (z_out_3(0)), (z_out_3(0)), STD_LOGIC_VECTOR'( QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_or_cse
      & and_dcpl_726 & and_937_ssc));
  QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_4_nl <= QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_3_nl
      AND nor_1324_seb;
  nor_1109_nl <= NOT((fsm_output(6)) OR mux_tmp_1440);
  nor_1110_nl <= NOT((NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT (fsm_output(2))));
  mux_1441_nl <= MUX_s_1_2_2(nor_1109_nl, nor_1110_nl, fsm_output(7));
  CACHE_UPDATE_LOOP_3_k_and_1_nl <= (NOT and_dcpl_629) AND mux_1441_nl AND and_dcpl_628;
  or_594_nl <= reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 OR reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  RMS_NORM_LOOP_2_2_mux1h_nl <= MUX1HOT_s_1_3_2(RMS_NORM_LOOP_2_2_unequal_tmp_mx0w0,
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1, or_594_nl, STD_LOGIC_VECTOR'(
      and_dcpl_386 & and_dcpl_629 & and_dcpl_207));
  nand_348_nl <= NOT((fsm_output(5)) AND and_1637_cse);
  or_2341_nl <= (NOT (fsm_output(5))) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(2));
  mux_1438_nl <= MUX_s_1_2_2(nand_348_nl, or_2341_nl, fsm_output(3));
  or_2342_nl <= (fsm_output(6)) OR mux_1438_nl;
  or_2340_nl <= (fsm_output(3)) OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (fsm_output(1))
      OR (fsm_output(2));
  or_2339_nl <= (fsm_output(3)) OR (NOT((fsm_output(5)) AND (fsm_output(2))));
  mux_1437_nl <= MUX_s_1_2_2(or_2340_nl, or_2339_nl, fsm_output(6));
  mux_1439_nl <= MUX_s_1_2_2(or_2342_nl, mux_1437_nl, fsm_output(7));
  RMS_NORM_LOOP_2_2_and_36_nl <= RMS_NORM_LOOP_2_2_mux1h_nl AND (NOT(mux_1439_nl
      OR or_tmp_48));
  GEMM_3D_FLOAT_LOOP_1_i_mux_1_nl <= MUX_s_1_2_2(RMS_NORM_LOOP_2_2_and_36_nl, (z_out_5(0)),
      GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c1);
  and_688_nl <= or_dcpl_1108 AND and_dcpl_202 AND and_dcpl_642;
  and_693_nl <= or_dcpl_1114 AND and_dcpl_202 AND and_dcpl_642;
  and_704_nl <= or_dcpl_1118 AND and_dcpl_202 AND and_dcpl_642;
  and_709_nl <= or_dcpl_1120 AND and_dcpl_202 AND and_dcpl_642;
  and_713_nl <= or_dcpl_1121 AND and_dcpl_202 AND and_dcpl_642;
  and_717_nl <= or_dcpl_1122 AND and_dcpl_202 AND and_dcpl_642;
  and_721_nl <= or_dcpl_1123 AND and_dcpl_202 AND and_dcpl_642;
  and_725_nl <= or_dcpl_1125 AND and_dcpl_202 AND and_dcpl_642;
  and_729_nl <= or_dcpl_1126 AND and_dcpl_202 AND and_dcpl_642;
  and_733_nl <= or_dcpl_1127 AND and_dcpl_202 AND and_dcpl_642;
  and_737_nl <= or_dcpl_1128 AND and_dcpl_202 AND and_dcpl_642;
  and_741_nl <= or_dcpl_1130 AND and_dcpl_202 AND and_dcpl_642;
  and_749_nl <= or_dcpl_1132 AND and_dcpl_202 AND and_dcpl_642;
  and_753_nl <= or_dcpl_1133 AND and_dcpl_202 AND and_dcpl_642;
  LINEAR_FORWARD_NO_MUL_LOOP_2_and_1_nl <= (LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1(4))
      AND LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4 AND (RMS_NORM_LOOP_2_2_i_4_0_sva_1(4));
  and_755_nl <= and_dcpl_215 AND nor_1138_m1c;
  nand_353_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 0)=STD_LOGIC_VECTOR'("1111111")));
  mux_1491_nl <= MUX_s_1_2_2(nand_353_nl, or_tmp_1218, fsm_output(7));
  nor_1136_nl <= NOT(mux_1491_nl OR (fsm_output(8)));
  and_757_nl <= and_dcpl_291 AND nor_1138_m1c;
  nand_356_nl <= NOT((fsm_output(5)) AND (fsm_output(0)) AND (fsm_output(2)) AND
      (NOT (fsm_output(4))));
  mux_1514_nl <= MUX_s_1_2_2((NOT and_1570_cse), or_tmp_1221, fsm_output(0));
  mux_1515_nl <= MUX_s_1_2_2(mux_1514_nl, mux_1513_cse, fsm_output(5));
  mux_1516_nl <= MUX_s_1_2_2(nand_356_nl, mux_1515_nl, fsm_output(3));
  nor_1141_nl <= NOT(RESHAPE_2D_TO_3D_LOOP_2_2_and_cse OR (fsm_output(3)) OR (NOT
      (fsm_output(4))) OR (fsm_output(6)));
  nor_1142_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(3))) OR (fsm_output(4))
      OR (NOT (fsm_output(6))));
  mux_1536_nl <= MUX_s_1_2_2(nor_1141_nl, nor_1142_nl, fsm_output(0));
  or_2463_nl <= (NOT (fsm_output(3))) OR (fsm_output(4)) OR (NOT (fsm_output(6)));
  or_2461_nl <= (z_out_4(2)) OR (fsm_output(3)) OR (NOT (fsm_output(4))) OR (fsm_output(6));
  mux_1534_nl <= MUX_s_1_2_2(or_2463_nl, or_2461_nl, fsm_output(1));
  nor_1143_nl <= NOT((fsm_output(0)) OR mux_1534_nl);
  mux_1537_nl <= MUX_s_1_2_2(mux_1536_nl, nor_1143_nl, fsm_output(2));
  APPLY_ROTARY_POS_EMB_LOOP_1_i_or_nl <= ((NOT mux_1309_cse) AND and_1559_cse AND
      nor_1026_cse AND and_dcpl_576) OR ((NOT mux_1516_nl) AND and_dcpl_718) OR (mux_1537_nl
      AND and_dcpl_388);
  APPLY_ROTARY_POS_EMB_LOOP_1_i_mux1h_5_nl <= MUX1HOT_s_1_5_2(and_28_cse, LINEAR_FORWARD_NO_MUL_LOOP_2_and_1_nl,
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1, RMS_NORM_LOOP_2_2_and_32_ssc_mx0w3,
      (z_out_4(0)), STD_LOGIC_VECTOR'( and_dcpl_363 & and_755_nl & nor_1136_nl &
      and_757_nl & APPLY_ROTARY_POS_EMB_LOOP_1_i_or_nl));
  attention_2_1_16_16_4_4_v_proj_re_mux1h_4_nl <= MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16_mx1,
      attention_2_1_16_16_4_4_v_proj_re_0_15_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_39_16,
      STD_LOGIC_VECTOR'( and_dcpl_725 & and_dcpl_726 & and_dcpl_410));
  not_4557_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_8_nl <= MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16_mx1,
      attention_2_1_16_16_4_4_v_proj_re_0_0_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_39_16,
      STD_LOGIC_VECTOR'( and_dcpl_725 & and_dcpl_726 & and_dcpl_410));
  not_4558_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_12_nl <= MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16_mx1,
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_39_16,
      STD_LOGIC_VECTOR'( and_dcpl_725 & and_dcpl_726 & and_dcpl_410));
  not_4559_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_16_nl <= MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16_mx1,
      attention_2_1_16_16_4_4_v_proj_re_0_3_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_39_16,
      STD_LOGIC_VECTOR'( and_dcpl_725 & and_dcpl_726 & and_dcpl_410));
  not_4560_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_20_nl <= MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16_mx1,
      attention_2_1_16_16_4_4_v_proj_re_0_7_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_39_16,
      STD_LOGIC_VECTOR'( and_dcpl_725 & and_dcpl_726 & and_dcpl_410));
  not_4561_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_21_nl <= MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16_mx1,
      attention_2_1_16_16_4_4_k_proj_re_0_7_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_7_sva_2_39_16,
      STD_LOGIC_VECTOR'( and_dcpl_725 & and_dcpl_726 & and_dcpl_410));
  not_4562_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_35_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_7_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_754);
  not_4441_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_34_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_8_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_760);
  not_4440_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_33_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_6_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_764);
  not_4439_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_32_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_9_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_768);
  not_4438_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_31_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_5_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_772);
  not_4437_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_30_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_10_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_776);
  not_4436_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_29_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_4_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_780);
  not_4435_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_28_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_11_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_784);
  not_4434_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_27_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_12_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_788);
  not_4433_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_26_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_13_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_792);
  not_4432_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_25_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_1_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_796);
  not_4431_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_24_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_14_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_800);
  not_4430_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_23_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_0_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_804);
  not_4429_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_22_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_15_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_812);
  not_4428_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_21_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_8_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_821);
  not_4427_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_20_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_6_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_827);
  not_4426_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_19_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_9_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_832);
  not_4425_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_18_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_5_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_837);
  not_4424_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_17_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_4_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_851);
  not_4422_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux_16_nl <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_15_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), and_dcpl_880);
  not_4415_nl <= NOT and_dcpl_619;
  and_1184_nl <= or_dcpl_1141 AND and_dcpl_191 AND and_dcpl_641 AND and_dcpl_813;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_40_nl <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_re_0_10_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16, STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16_mx0c1
      & and_dcpl_843 & and_dcpl_207 & and_dcpl_847));
  not_4423_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_42_nl <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_re_0_11_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16, STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16_mx0c1
      & and_dcpl_856 & and_dcpl_207 & and_dcpl_847));
  not_4421_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_43_nl <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_re_0_12_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16, STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16_mx0c1
      & and_dcpl_860 & and_dcpl_207 & and_dcpl_847));
  not_4420_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_44_nl <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_re_0_13_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16, STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16_mx0c1
      & and_dcpl_864 & and_dcpl_207 & and_dcpl_847));
  not_4419_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_45_nl <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_re_0_1_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16, STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16_mx0c1
      & and_dcpl_868 & and_dcpl_207 & and_dcpl_847));
  not_4418_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_46_nl <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_re_0_14_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16, STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16_mx0c1
      & and_dcpl_872 & and_dcpl_207 & and_dcpl_847));
  not_4417_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_47_nl <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_re_0_0_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16, STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16_mx0c1
      & and_dcpl_876 & and_dcpl_207 & and_dcpl_847));
  not_4416_nl <= NOT and_dcpl_619;
  GEMM_3D_FLOAT_LOOP_4_l_GEMM_3D_FLOAT_LOOP_4_l_mux_nl <= MUX_s_1_2_2((z_out_5(1)),
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0)), APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c2);
  RMS_NORM_LOOP_2_2_mux_23_nl <= MUX_s_1_16_2('1', '0', '1', '1', '1', '1', '1',
      '1', '1', '1', '1', '1', '1', '1', '1', '1', reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
      & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  and_1810_nl <= or_1907_cse AND (fsm_output(4));
  mux_2242_nl <= MUX_s_1_2_2(nor_tmp_289, and_1810_nl, fsm_output(0));
  mux_2243_nl <= MUX_s_1_2_2((NOT mux_2242_nl), nor_tmp_329, fsm_output(5));
  mux_2244_nl <= MUX_s_1_2_2((NOT (fsm_output(5))), mux_2243_nl, fsm_output(3));
  mux_2245_nl <= MUX_s_1_2_2(mux_2244_nl, mux_tmp_1027, or_3039_cse);
  and_1254_nl <= (NOT mux_2245_nl) AND and_dcpl_413;
  RMS_NORM_LOOP_1_1_mux1h_nl <= MUX1HOT_s_1_3_2(RMS_NORM_LOOP_2_2_mux_23_nl, reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1,
      (NOT QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1), STD_LOGIC_VECTOR'(
      and_dcpl_448 & and_1254_nl & and_dcpl_557));
  nor_1316_nl <= NOT((fsm_output(5)) OR (or_1732_cse AND CONV_SL_1_1(fsm_output(4
      DOWNTO 3)=STD_LOGIC_VECTOR'("11"))));
  and_1809_nl <= (fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(3)) AND (fsm_output(4));
  mux_2239_nl <= MUX_s_1_2_2(nand_381_cse, and_1809_nl, fsm_output(5));
  mux_2240_nl <= MUX_s_1_2_2(nor_1316_nl, mux_2239_nl, fsm_output(2));
  nor_1320_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(6)) OR mux_2240_nl);
  or_3033_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"));
  or_3032_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"));
  mux_2238_nl <= MUX_s_1_2_2(or_3033_nl, or_3032_nl, fsm_output(6));
  nor_1321_nl <= NOT((fsm_output(8)) OR mux_2238_nl);
  mux_2241_nl <= MUX_s_1_2_2(nor_1320_nl, nor_1321_nl, fsm_output(7));
  RMS_NORM_LOOP_1_1_or_nl <= (RMS_NORM_LOOP_1_1_mux1h_nl AND mux_2241_nl) OR (and_dcpl_241
      AND and_dcpl_293);
  GEMM_3D_FLOAT_LOOP_4_l_or_1_nl <= and_dcpl_726 OR APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c4;
  GEMM_3D_FLOAT_LOOP_4_l_mux1h_13_nl <= MUX1HOT_s_1_3_2((z_out_5(0)), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2,
      RMS_NORM_LOOP_1_1_or_nl, STD_LOGIC_VECTOR'( GEMM_3D_FLOAT_LOOP_4_l_or_1_nl
      & APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c2 & APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c3));
  and_939_nl <= and_dcpl_732 AND and_dcpl_875;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_26_nl <= MUX1HOT_v_16_4_2(z_out_1, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0,
      STD_LOGIC_VECTOR'( and_939_nl & and_dcpl_876 & and_dcpl_207 & and_dcpl_847));
  not_4471_nl <= NOT and_dcpl_619;
  or_3191_nl <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(0))) OR mux_1639_cse;
  mux_1640_nl <= MUX_s_1_2_2(or_2699_cse, or_3191_nl, and_1773_cse);
  or_3192_nl <= (fsm_output(7)) OR (NOT mux_1640_nl);
  mux_1641_nl <= MUX_s_1_2_2(nand_365_cse, or_3192_nl, fsm_output(6));
  and_941_nl <= and_dcpl_732 AND and_dcpl_867;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_28_nl <= MUX1HOT_v_16_4_2(z_out_1, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0,
      STD_LOGIC_VECTOR'( and_941_nl & and_dcpl_868 & and_dcpl_207 & and_dcpl_847));
  not_4470_nl <= NOT and_dcpl_619;
  or_3194_nl <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(0))) OR mux_1639_cse;
  mux_1643_nl <= MUX_s_1_2_2(or_2699_cse, or_3194_nl, and_1773_cse);
  or_3195_nl <= (fsm_output(7)) OR (NOT mux_1643_nl);
  mux_1644_nl <= MUX_s_1_2_2(nand_365_cse, or_3195_nl, fsm_output(6));
  and_958_nl <= and_dcpl_732 AND and_dcpl_879;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_40_nl <= MUX1HOT_v_16_4_2(z_out_1, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0,
      STD_LOGIC_VECTOR'( and_958_nl & and_dcpl_880 & and_dcpl_207 & and_dcpl_847));
  not_4464_nl <= NOT and_dcpl_619;
  nand_81_nl <= NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      AND CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(0)) AND (NOT mux_1639_cse));
  mux_1726_nl <= MUX_s_1_2_2(or_2699_cse, nand_81_nl, and_1773_cse);
  or_3197_nl <= (fsm_output(7)) OR (NOT mux_1726_nl);
  mux_1727_nl <= MUX_s_1_2_2(nand_365_cse, or_3197_nl, fsm_output(6));
  attention_2_1_16_16_4_4_k_proj_re_mux_43_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_804);
  not_4458_nl <= NOT and_dcpl_619;
  or_2491_nl <= reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 OR CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd/=STD_LOGIC_VECTOR'("000"));
  mux_1813_nl <= MUX_s_1_2_2(mux_1812_cse, mux_806_cse, or_2491_nl);
  mux_1814_nl <= MUX_s_1_2_2(or_2249_cse, mux_1813_nl, and_1773_cse);
  mux_1815_nl <= MUX_s_1_2_2(mux_1814_nl, mux_1809_cse, fsm_output(4));
  mux_1816_nl <= MUX_s_1_2_2(mux_1815_nl, or_1983_cse, fsm_output(5));
  attention_2_1_16_16_4_4_k_proj_re_mux_42_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_796);
  not_4457_nl <= NOT and_dcpl_619;
  or_2490_nl <= (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) OR CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd/=STD_LOGIC_VECTOR'("000"));
  mux_1822_nl <= MUX_s_1_2_2(mux_1812_cse, mux_806_cse, or_2490_nl);
  mux_1823_nl <= MUX_s_1_2_2(or_2249_cse, mux_1822_nl, and_1773_cse);
  mux_1824_nl <= MUX_s_1_2_2(mux_1823_nl, mux_1809_cse, fsm_output(4));
  mux_1825_nl <= MUX_s_1_2_2(mux_1824_nl, or_1983_cse, fsm_output(5));
  attention_2_1_16_16_4_4_k_proj_re_mux_41_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_776);
  not_4456_nl <= NOT and_dcpl_619;
  nor_514_nl <= NOT(CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)/=STD_LOGIC_VECTOR'("10")) OR reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 OR
      (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0))));
  mux_1831_nl <= MUX_s_1_2_2(mux_806_cse, mux_1812_cse, nor_514_nl);
  mux_1832_nl <= MUX_s_1_2_2(or_2249_cse, mux_1831_nl, and_1773_cse);
  mux_1833_nl <= MUX_s_1_2_2(mux_1832_nl, mux_1809_cse, fsm_output(4));
  mux_1834_nl <= MUX_s_1_2_2(mux_1833_nl, or_1983_cse, fsm_output(5));
  attention_2_1_16_16_4_4_k_proj_re_mux_40_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_784);
  not_4455_nl <= NOT and_dcpl_619;
  and_1727_nl <= CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"))
      AND reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 AND (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0));
  mux_1840_nl <= MUX_s_1_2_2(mux_806_cse, mux_1812_cse, and_1727_nl);
  mux_1841_nl <= MUX_s_1_2_2(or_2249_cse, mux_1840_nl, and_1773_cse);
  mux_1842_nl <= MUX_s_1_2_2(mux_1841_nl, mux_1809_cse, fsm_output(4));
  mux_1843_nl <= MUX_s_1_2_2(mux_1842_nl, or_1983_cse, fsm_output(5));
  attention_2_1_16_16_4_4_k_proj_re_mux_39_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_788);
  not_4454_nl <= NOT and_dcpl_619;
  or_2653_nl <= CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("11"))
      OR reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 OR (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0));
  mux_1849_nl <= MUX_s_1_2_2(mux_1812_cse, mux_806_cse, or_2653_nl);
  mux_1850_nl <= MUX_s_1_2_2(or_2249_cse, mux_1849_nl, and_1773_cse);
  mux_1851_nl <= MUX_s_1_2_2(mux_1850_nl, mux_1809_cse, fsm_output(4));
  mux_1852_nl <= MUX_s_1_2_2(mux_1851_nl, or_1983_cse, fsm_output(5));
  attention_2_1_16_16_4_4_k_proj_re_mux_38_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_792);
  not_4453_nl <= NOT and_dcpl_619;
  nand_369_nl <= NOT(CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)=STD_LOGIC_VECTOR'("11")) AND reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 AND
      (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0))));
  mux_1858_nl <= MUX_s_1_2_2(mux_1812_cse, mux_806_cse, nand_369_nl);
  mux_1859_nl <= MUX_s_1_2_2(or_2249_cse, mux_1858_nl, and_1773_cse);
  mux_1860_nl <= MUX_s_1_2_2(mux_1859_nl, mux_1809_cse, fsm_output(4));
  mux_1861_nl <= MUX_s_1_2_2(mux_1860_nl, or_1983_cse, fsm_output(5));
  attention_2_1_16_16_4_4_k_proj_re_mux_37_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_800);
  not_4452_nl <= NOT and_dcpl_619;
  and_1658_nl <= (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) AND CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd=STD_LOGIC_VECTOR'("111"));
  mux_1867_nl <= MUX_s_1_2_2(mux_806_cse, mux_1812_cse, and_1658_nl);
  mux_1868_nl <= MUX_s_1_2_2(or_2249_cse, mux_1867_nl, and_1773_cse);
  mux_1869_nl <= MUX_s_1_2_2(mux_1868_nl, mux_1809_cse, fsm_output(4));
  mux_1870_nl <= MUX_s_1_2_2(mux_1869_nl, or_1983_cse, fsm_output(5));
  attention_2_1_16_16_4_4_k_proj_re_mux_36_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_812);
  not_4451_nl <= NOT and_dcpl_619;
  and_1733_nl <= CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
      AND reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 AND (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0))
      AND (fsm_output(0));
  mux_1874_nl <= MUX_s_1_2_2(mux_806_cse, or_2249_cse, and_1733_nl);
  or_2664_nl <= (NOT (LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1(4))) OR (fsm_output(0));
  mux_1873_nl <= MUX_s_1_2_2(or_1983_cse, mux_806_cse, or_2664_nl);
  mux_1875_nl <= MUX_s_1_2_2(mux_1874_nl, mux_1873_nl, fsm_output(1));
  mux_1876_nl <= MUX_s_1_2_2(or_2249_cse, mux_1875_nl, and_1773_cse);
  mux_1877_nl <= MUX_s_1_2_2(mux_1876_nl, mux_1809_cse, fsm_output(4));
  mux_1878_nl <= MUX_s_1_2_2(mux_1877_nl, or_1983_cse, fsm_output(5));
  attention_2_1_16_16_4_4_k_proj_re_mux_35_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_959);
  not_4450_nl <= NOT and_dcpl_619;
  nor_524_nl <= NOT(CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)/=STD_LOGIC_VECTOR'("00")) OR (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1)
      OR (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0))));
  mux_1884_nl <= MUX_s_1_2_2(mux_806_cse, mux_1812_cse, nor_524_nl);
  mux_1885_nl <= MUX_s_1_2_2(or_2249_cse, mux_1884_nl, and_1773_cse);
  mux_1886_nl <= MUX_s_1_2_2(mux_1885_nl, mux_1809_cse, fsm_output(4));
  mux_1887_nl <= MUX_s_1_2_2(mux_1886_nl, or_1983_cse, fsm_output(5));
  attention_2_1_16_16_4_4_k_proj_re_mux_34_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_780);
  not_4449_nl <= NOT and_dcpl_619;
  mux_1893_nl <= MUX_s_1_2_2(mux_1812_cse, mux_806_cse, or_2671_cse);
  mux_1894_nl <= MUX_s_1_2_2(or_2249_cse, mux_1893_nl, and_1773_cse);
  mux_1895_nl <= MUX_s_1_2_2(mux_1894_nl, mux_1809_cse, fsm_output(4));
  mux_1896_nl <= MUX_s_1_2_2(mux_1895_nl, or_1983_cse, fsm_output(5));
  attention_2_1_16_16_4_4_k_proj_re_mux_33_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_772);
  not_4448_nl <= NOT and_dcpl_619;
  or_2675_nl <= CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) OR (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0));
  mux_1902_nl <= MUX_s_1_2_2(mux_1812_cse, mux_806_cse, or_2675_nl);
  mux_1903_nl <= MUX_s_1_2_2(or_2249_cse, mux_1902_nl, and_1773_cse);
  mux_1904_nl <= MUX_s_1_2_2(mux_1903_nl, mux_1809_cse, fsm_output(4));
  mux_1905_nl <= MUX_s_1_2_2(mux_1904_nl, or_1983_cse, fsm_output(5));
  attention_2_1_16_16_4_4_k_proj_re_mux_32_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_764);
  not_4447_nl <= NOT and_dcpl_619;
  nor_441_nl <= NOT(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 OR CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd/=STD_LOGIC_VECTOR'("011")));
  mux_1911_nl <= MUX_s_1_2_2(mux_806_cse, mux_1812_cse, nor_441_nl);
  mux_1912_nl <= MUX_s_1_2_2(or_2249_cse, mux_1911_nl, and_1773_cse);
  mux_1913_nl <= MUX_s_1_2_2(mux_1912_nl, mux_1809_cse, fsm_output(4));
  mux_1914_nl <= MUX_s_1_2_2(mux_1913_nl, or_1983_cse, fsm_output(5));
  attention_2_1_16_16_4_4_k_proj_re_mux_31_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_754);
  not_4446_nl <= NOT and_dcpl_619;
  and_1656_nl <= reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 AND CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd=STD_LOGIC_VECTOR'("011"));
  mux_1920_nl <= MUX_s_1_2_2(mux_806_cse, mux_1812_cse, and_1656_nl);
  mux_1921_nl <= MUX_s_1_2_2(or_2249_cse, mux_1920_nl, and_1773_cse);
  mux_1922_nl <= MUX_s_1_2_2(mux_1921_nl, mux_1809_cse, fsm_output(4));
  mux_1923_nl <= MUX_s_1_2_2(mux_1922_nl, or_1983_cse, fsm_output(5));
  attention_2_1_16_16_4_4_k_proj_re_mux_30_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_760);
  not_4445_nl <= NOT and_dcpl_619;
  mux_1929_nl <= MUX_s_1_2_2(mux_1812_cse, mux_806_cse, or_2486_cse);
  mux_1930_nl <= MUX_s_1_2_2(or_2249_cse, mux_1929_nl, and_1773_cse);
  mux_1931_nl <= MUX_s_1_2_2(mux_1930_nl, mux_1809_cse, fsm_output(4));
  mux_1932_nl <= MUX_s_1_2_2(mux_1931_nl, or_1983_cse, fsm_output(5));
  attention_2_1_16_16_4_4_k_proj_re_mux_29_nl <= MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg(15
      DOWNTO 0)), and_dcpl_768);
  not_4444_nl <= NOT and_dcpl_619;
  or_2487_nl <= (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) OR CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd/=STD_LOGIC_VECTOR'("100"));
  mux_1938_nl <= MUX_s_1_2_2(mux_1812_cse, mux_806_cse, or_2487_nl);
  mux_1939_nl <= MUX_s_1_2_2(or_2249_cse, mux_1938_nl, and_1773_cse);
  mux_1940_nl <= MUX_s_1_2_2(mux_1939_nl, mux_1809_cse, fsm_output(4));
  mux_1941_nl <= MUX_s_1_2_2(mux_1940_nl, or_1983_cse, fsm_output(5));
  and_1025_nl <= and_dcpl_732 AND and_dcpl_585 AND and_dcpl_335;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_66_nl <= MUX1HOT_v_16_4_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_15_0, attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0, STD_LOGIC_VECTOR'( and_1025_nl
      & and_dcpl_983 & and_dcpl_240 & and_dcpl_626));
  not_4563_nl <= NOT and_dcpl_619;
  nor_533_nl <= NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1/=STD_LOGIC_VECTOR'("00"))
      OR (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd));
  mux_1946_nl <= MUX_s_1_2_2(mux_tmp_1945, mux_tmp_1943, nor_533_nl);
  and_1031_nl <= and_dcpl_732 AND and_dcpl_585 AND and_dcpl_480;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_67_nl <= MUX1HOT_v_16_4_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_15_0, attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0, STD_LOGIC_VECTOR'( and_1031_nl
      & and_dcpl_983 & and_dcpl_240 & and_dcpl_626));
  not_4564_nl <= NOT and_dcpl_619;
  nor_535_nl <= NOT((NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2)
      OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1/=STD_LOGIC_VECTOR'("00"))
      OR (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd));
  mux_1947_nl <= MUX_s_1_2_2(mux_tmp_1945, mux_tmp_1943, nor_535_nl);
  attention_2_1_16_16_4_4_k_proj_re_mux1h_69_nl <= MUX1HOT_v_8_7_2((drf_output_sdt_2_sva_15_0_mx0w0(15
      DOWNTO 8)), (attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_15_0(15 DOWNTO 8)),
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0_mx0w1(15 DOWNTO 8)), (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(15
      DOWNTO 8)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8,
      (output_0_3_lpi_3_15_0(15 DOWNTO 8)), (drf_output_sdt_3_sva_15_0_mx0w3(15 DOWNTO
      8)), STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c1
      & and_dcpl_983 & and_dcpl_240 & and_dcpl_626 & and_dcpl_207 & and_dcpl_739
      & apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c8));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_119_nl <= MUX1HOT_v_8_7_2((drf_output_sdt_2_sva_15_0_mx0w0(7
      DOWNTO 0)), (attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_15_0(7 DOWNTO 0)),
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0_mx0w1(7 DOWNTO 0)), (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(7
      DOWNTO 0)), STD_LOGIC_VECTOR'( APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7
      & APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6
      & APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5
      & APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4
      & APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3
      & APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2
      & APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1
      & APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0),
      (output_0_3_lpi_3_15_0(7 DOWNTO 0)), (drf_output_sdt_3_sva_15_0_mx0w3(7 DOWNTO
      0)), STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c1
      & and_dcpl_983 & and_dcpl_240 & and_dcpl_626 & and_dcpl_207 & and_dcpl_739
      & apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c8));
  not_4565_nl <= NOT and_dcpl_619;
  nor_1203_nl <= NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(7))) OR (fsm_output(8)));
  nor_1204_nl <= NOT(and_1474_cse OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01")));
  mux_1970_nl <= MUX_s_1_2_2(nor_1203_nl, nor_1204_nl, fsm_output(2));
  nor_1201_nl <= NOT((NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd OR
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("11"))))
      OR (NOT (fsm_output(0))) OR (fsm_output(7)) OR (NOT (fsm_output(8))));
  nor_1202_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10")));
  mux_1969_nl <= MUX_s_1_2_2(nor_1201_nl, nor_1202_nl, fsm_output(1));
  and_1749_nl <= (fsm_output(2)) AND mux_1969_nl;
  mux_1971_nl <= MUX_s_1_2_2(mux_1970_nl, and_1749_nl, fsm_output(3));
  and_1753_nl <= (fsm_output(4)) AND mux_1971_nl;
  nor_1206_nl <= NOT((CONV_SL_1_1(fsm_output(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1111")))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10")));
  mux_1972_nl <= MUX_s_1_2_2(and_1753_nl, nor_1206_nl, fsm_output(5));
  and_1754_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11")) AND
      (NOT((NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd OR (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1))
      OR (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2) OR (NOT (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0)))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")))) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))));
  mux_1967_nl <= MUX_s_1_2_2(and_1754_nl, and_dcpl_26, fsm_output(4));
  nor_1208_nl <= NOT((fsm_output(4)) OR and_1638_cse OR CONV_SL_1_1(fsm_output(8
      DOWNTO 7)/=STD_LOGIC_VECTOR'("00")));
  mux_1968_nl <= MUX_s_1_2_2(mux_1967_nl, nor_1208_nl, fsm_output(5));
  mux_1973_nl <= MUX_s_1_2_2(mux_1972_nl, mux_1968_nl, fsm_output(6));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_70_nl <= MUX1HOT_v_8_3_2((z_out(15 DOWNTO
      8)), (rms_norm_16_div_cmp_z_oreg(15 DOWNTO 8)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm,
      STD_LOGIC_VECTOR'( and_1042_ssc & and_dcpl_999 & and_dcpl_374));
  not_5074_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_128_nl <= MUX1HOT_s_1_3_2((z_out(7)), (rms_norm_16_div_cmp_z_oreg(7)),
      APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm,
      STD_LOGIC_VECTOR'( and_1042_ssc & and_dcpl_999 & and_dcpl_374));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_129_nl <= MUX1HOT_s_1_3_2((z_out(6)), (rms_norm_16_div_cmp_z_oreg(6)),
      APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm,
      STD_LOGIC_VECTOR'( and_1042_ssc & and_dcpl_999 & and_dcpl_374));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_130_nl <= MUX1HOT_s_1_3_2((z_out(5)), (rms_norm_16_div_cmp_z_oreg(5)),
      APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm,
      STD_LOGIC_VECTOR'( and_1042_ssc & and_dcpl_999 & and_dcpl_374));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_131_nl <= MUX1HOT_s_1_3_2((z_out(4)), (rms_norm_16_div_cmp_z_oreg(4)),
      APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm,
      STD_LOGIC_VECTOR'( and_1042_ssc & and_dcpl_999 & and_dcpl_374));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_132_nl <= MUX1HOT_s_1_3_2((z_out(3)), (rms_norm_16_div_cmp_z_oreg(3)),
      APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm,
      STD_LOGIC_VECTOR'( and_1042_ssc & and_dcpl_999 & and_dcpl_374));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_133_nl <= MUX1HOT_s_1_3_2((z_out(2)), (rms_norm_16_div_cmp_z_oreg(2)),
      APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm,
      STD_LOGIC_VECTOR'( and_1042_ssc & and_dcpl_999 & and_dcpl_374));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_134_nl <= MUX1HOT_s_1_3_2((z_out(1)), (rms_norm_16_div_cmp_z_oreg(1)),
      APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm,
      STD_LOGIC_VECTOR'( and_1042_ssc & and_dcpl_999 & and_dcpl_374));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_135_nl <= MUX1HOT_s_1_3_2((z_out(0)), (rms_norm_16_div_cmp_z_oreg(0)),
      APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm,
      STD_LOGIC_VECTOR'( and_1042_ssc & and_dcpl_999 & and_dcpl_374));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_71_nl <= MUX1HOT_v_8_3_2((z_out_1(15 DOWNTO
      8)), (rms_norm_16_div_cmp_z_oreg(15 DOWNTO 8)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm,
      STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1
      & and_dcpl_1003 & and_dcpl_207));
  not_5066_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_120_nl <= MUX1HOT_s_1_3_2((z_out_1(7)),
      (rms_norm_16_div_cmp_z_oreg(7)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm,
      STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1
      & and_dcpl_1003 & and_dcpl_207));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_121_nl <= MUX1HOT_s_1_3_2((z_out_1(6)),
      (rms_norm_16_div_cmp_z_oreg(6)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm,
      STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1
      & and_dcpl_1003 & and_dcpl_207));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_122_nl <= MUX1HOT_s_1_3_2((z_out_1(5)),
      (rms_norm_16_div_cmp_z_oreg(5)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm,
      STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1
      & and_dcpl_1003 & and_dcpl_207));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_123_nl <= MUX1HOT_s_1_3_2((z_out_1(4)),
      (rms_norm_16_div_cmp_z_oreg(4)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm,
      STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1
      & and_dcpl_1003 & and_dcpl_207));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_124_nl <= MUX1HOT_s_1_3_2((z_out_1(3)),
      (rms_norm_16_div_cmp_z_oreg(3)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm,
      STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1
      & and_dcpl_1003 & and_dcpl_207));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_125_nl <= MUX1HOT_s_1_3_2((z_out_1(2)),
      (rms_norm_16_div_cmp_z_oreg(2)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm,
      STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1
      & and_dcpl_1003 & and_dcpl_207));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_126_nl <= MUX1HOT_s_1_3_2((z_out_1(1)),
      (rms_norm_16_div_cmp_z_oreg(1)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm,
      STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1
      & and_dcpl_1003 & and_dcpl_207));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_127_nl <= MUX1HOT_s_1_3_2((z_out_1(0)),
      (rms_norm_16_div_cmp_z_oreg(0)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm,
      STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1
      & and_dcpl_1003 & and_dcpl_207));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_72_nl <= MUX1HOT_v_16_5_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_15_0, z_out_1, output_0_0_lpi_3_15_0,
      drf_output_sdt_3_sva_15_0_mx0w3, STD_LOGIC_VECTOR'( attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c1
      & and_dcpl_410 & and_dcpl_240 & and_dcpl_739 & attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c6));
  not_4566_nl <= NOT and_dcpl_619;
  mux_2010_nl <= MUX_s_1_2_2(mux_304_cse, or_2457_cse, fsm_output(3));
  nand_93_nl <= NOT((fsm_output(4)) AND (NOT mux_2010_nl));
  mux_2009_nl <= MUX_s_1_2_2(mux_tmp_919, or_1197_cse, fsm_output(4));
  mux_2011_nl <= MUX_s_1_2_2(nand_93_nl, mux_2009_nl, fsm_output(5));
  nand_92_nl <= NOT((fsm_output(3)) AND (NOT((NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd
      OR (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1)) OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2
      OR (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0)) OR CONV_SL_1_1(fsm_output(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")))) OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")))));
  mux_2005_nl <= MUX_s_1_2_2(mux_304_cse, or_2457_cse, and_1474_cse);
  and_1759_nl <= or_3039_cse AND (fsm_output(0));
  mux_2002_nl <= MUX_s_1_2_2(or_2457_cse, mux_tmp_919, and_1759_nl);
  mux_2003_nl <= MUX_s_1_2_2(mux_2002_nl, mux_tmp_919, fsm_output(1));
  mux_2006_nl <= MUX_s_1_2_2(mux_2005_nl, mux_2003_nl, fsm_output(3));
  mux_2007_nl <= MUX_s_1_2_2(nand_92_nl, mux_2006_nl, fsm_output(4));
  mux_2000_nl <= MUX_s_1_2_2(mux_tmp_919, or_1197_cse, and_dcpl_65);
  or_2720_nl <= and_dcpl_65 OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100"));
  mux_2001_nl <= MUX_s_1_2_2(mux_2000_nl, or_2720_nl, fsm_output(4));
  mux_2008_nl <= MUX_s_1_2_2(mux_2007_nl, mux_2001_nl, fsm_output(5));
  mux_2012_nl <= MUX_s_1_2_2(mux_2011_nl, mux_2008_nl, fsm_output(2));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_73_nl <= MUX1HOT_v_16_3_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_15_0, z_out, STD_LOGIC_VECTOR'(
      attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0_mx0c1 & and_dcpl_410 & and_dcpl_240));
  not_4567_nl <= NOT and_dcpl_619;
  mux_2021_nl <= MUX_s_1_2_2(mux_tmp_2015, mux_tmp_2013, fsm_output(3));
  or_2733_nl <= and_1762_cse OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  and_1763_nl <= (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd) AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1))
      AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0))
      AND (fsm_output(0));
  mux_2018_nl <= MUX_s_1_2_2(or_2733_nl, mux_tmp_2013, and_1763_nl);
  mux_2019_nl <= MUX_s_1_2_2(mux_tmp_2015, mux_2018_nl, fsm_output(3));
  mux_2016_nl <= MUX_s_1_2_2(mux_tmp_2015, mux_tmp_2013, fsm_output(0));
  mux_2017_nl <= MUX_s_1_2_2(mux_2016_nl, or_tmp_914, fsm_output(3));
  mux_2020_nl <= MUX_s_1_2_2(mux_2019_nl, mux_2017_nl, fsm_output(1));
  mux_2022_nl <= MUX_s_1_2_2(mux_2021_nl, mux_2020_nl, fsm_output(2));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_nl <= MUX_v_8_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(15
      DOWNTO 8)), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(15 DOWNTO 8)), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0(15
      DOWNTO 8)), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0(15 DOWNTO
      8)), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3(15 DOWNTO 8)), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm(15
      DOWNTO 8)), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_15_8, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_8,
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3(15 DOWNTO 8)), (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm(15
      DOWNTO 8)), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_15_8, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_8,
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3(15 DOWNTO 8)), (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm(15
      DOWNTO 8)), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_15_8, reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_ftd,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_74_nl <= MUX1HOT_v_8_9_2((drf_output_sdt_2_sva_15_0_mx0w0(15
      DOWNTO 8)), reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_ftd, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_15_8,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_15_8, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_ftd, APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_nl,
      output_0_1_lpi_3_15_8, (drf_output_sdt_3_sva_15_0_mx0w3(15 DOWNTO 8)), STD_LOGIC_VECTOR'(
      and_1055_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847 & and_dcpl_583 & and_dcpl_739 & and_1059_ssc));
  not_5054_nl <= NOT and_dcpl_619;
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_67_nl <= MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(7)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(7)), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0(7)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0(7)), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3(7)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm(7)), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_7,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_7, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3(7)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm(7)), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_7,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3(7)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm(7)), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_7,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_117_nl <= MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0(7)),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_7,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_7, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd, APPLY_ROTARY_POS_EMB_LOOP_6_mux_67_nl,
      output_0_1_lpi_3_7, (drf_output_sdt_3_sva_15_0_mx0w3(7)), STD_LOGIC_VECTOR'(
      and_1055_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847 & and_dcpl_583 & and_dcpl_739 & and_1059_ssc));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_88_nl <= MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(6)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(6)), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0(6)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0(6)), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3(6)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm(6)), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_6,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_6, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3(6)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm(6)), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_6,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_1, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3(6)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm(6)), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_6,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_1, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_152_nl <= MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0(6)),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_1, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_6,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_6, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_1, APPLY_ROTARY_POS_EMB_LOOP_6_mux_88_nl,
      output_0_1_lpi_3_6, (drf_output_sdt_3_sva_15_0_mx0w3(6)), STD_LOGIC_VECTOR'(
      and_1055_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847 & and_dcpl_583 & and_dcpl_739 & and_1059_ssc));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_89_nl <= MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(5)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(5)), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0(5)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0(5)), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3(5)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm(5)), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_5,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_5, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3(5)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm(5)), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_5,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_2, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3(5)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm(5)), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_5,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_2, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_153_nl <= MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0(5)),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_2, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_5,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_5, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_2, APPLY_ROTARY_POS_EMB_LOOP_6_mux_89_nl,
      output_0_1_lpi_3_5, (drf_output_sdt_3_sva_15_0_mx0w3(5)), STD_LOGIC_VECTOR'(
      and_1055_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847 & and_dcpl_583 & and_dcpl_739 & and_1059_ssc));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_90_nl <= MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(4)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(4)), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0(4)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0(4)), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3(4)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm(4)), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_4,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_4, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3(4)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm(4)), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_4,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_3, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3(4)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm(4)), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_4,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_3, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_154_nl <= MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0(4)),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_3, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_4,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_4, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_3, APPLY_ROTARY_POS_EMB_LOOP_6_mux_90_nl,
      output_0_1_lpi_3_4, (drf_output_sdt_3_sva_15_0_mx0w3(4)), STD_LOGIC_VECTOR'(
      and_1055_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847 & and_dcpl_583 & and_dcpl_739 & and_1059_ssc));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_91_nl <= MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(3)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(3)), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0(3)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0(3)), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3(3)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm(3)), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_3,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_3, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3(3)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm(3)), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_3,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_4, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3(3)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm(3)), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_3,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_4, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_155_nl <= MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0(3)),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_4, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_3,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_3, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_4, APPLY_ROTARY_POS_EMB_LOOP_6_mux_91_nl,
      output_0_1_lpi_3_3, (drf_output_sdt_3_sva_15_0_mx0w3(3)), STD_LOGIC_VECTOR'(
      and_1055_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847 & and_dcpl_583 & and_dcpl_739 & and_1059_ssc));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_92_nl <= MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(2)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(2)), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0(2)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0(2)), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3(2)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm(2)), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_2,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_2, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3(2)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm(2)), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_2,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_5, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3(2)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm(2)), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_2,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_5, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_156_nl <= MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0(2)),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_5, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_2,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_2, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_5, APPLY_ROTARY_POS_EMB_LOOP_6_mux_92_nl,
      output_0_1_lpi_3_2, (drf_output_sdt_3_sva_15_0_mx0w3(2)), STD_LOGIC_VECTOR'(
      and_1055_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847 & and_dcpl_583 & and_dcpl_739 & and_1059_ssc));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_93_nl <= MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(1)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(1)), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0(1)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0(1)), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3(1)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm(1)), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_1, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3(1)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm(1)), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_1,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_6, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3(1)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm(1)), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_1,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_6, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_157_nl <= MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0(1)),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_6, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_1,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_1, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_6, APPLY_ROTARY_POS_EMB_LOOP_6_mux_93_nl,
      output_0_1_lpi_3_1, (drf_output_sdt_3_sva_15_0_mx0w3(1)), STD_LOGIC_VECTOR'(
      and_1055_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847 & and_dcpl_583 & and_dcpl_739 & and_1059_ssc));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_94_nl <= MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1(0)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(0)), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0(0)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0(0)), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3(0)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm(0)), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_0,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_0, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3(0)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm(0)), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_0,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_7, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3(0)),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm(0)), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_0,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_7, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_158_nl <= MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0(0)),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_7, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_0,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_0, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_7, APPLY_ROTARY_POS_EMB_LOOP_6_mux_94_nl,
      output_0_1_lpi_3_0, (drf_output_sdt_3_sva_15_0_mx0w3(0)), STD_LOGIC_VECTOR'(
      and_1055_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847 & and_dcpl_583 & and_dcpl_739 & and_1059_ssc));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_75_nl <= MUX1HOT_v_3_6_2((drf_output_sdt_2_sva_15_0_mx0w0(15
      DOWNTO 13)), attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_13, attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_15_13,
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_15_13, apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_13,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_13, STD_LOGIC_VECTOR'(
      and_1060_itm & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847));
  not_4569_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_116_nl <= MUX1HOT_v_5_7_2((drf_output_sdt_2_sva_15_0_mx0w0(12
      DOWNTO 8)), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(12 DOWNTO 8)),
      (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0(12 DOWNTO 8)), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0(12
      DOWNTO 8)), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_12_8,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_12_8, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm(12
      DOWNTO 8)), STD_LOGIC_VECTOR'( and_1060_itm & and_dcpl_1011 & and_dcpl_983
      & and_dcpl_240 & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_144_nl <= MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0(7)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(7)), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0(7)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0(7)), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_7, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm(7)),
      STD_LOGIC_VECTOR'( and_1060_itm & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240
      & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_145_nl <= MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0(6)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(6)), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0(6)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0(6)), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_6, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm(6)),
      STD_LOGIC_VECTOR'( and_1060_itm & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240
      & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_146_nl <= MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0(5)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(5)), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0(5)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0(5)), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_5, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm(5)),
      STD_LOGIC_VECTOR'( and_1060_itm & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240
      & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_147_nl <= MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0(4)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(4)), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0(4)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0(4)), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_4, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm(4)),
      STD_LOGIC_VECTOR'( and_1060_itm & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240
      & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_148_nl <= MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0(3)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(3)), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0(3)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0(3)), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_3, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm(3)),
      STD_LOGIC_VECTOR'( and_1060_itm & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240
      & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_149_nl <= MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0(2)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(2)), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0(2)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0(2)), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_2, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm(2)),
      STD_LOGIC_VECTOR'( and_1060_itm & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240
      & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_150_nl <= MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0(1)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(1)), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0(1)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0(1)), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_1, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm(1)),
      STD_LOGIC_VECTOR'( and_1060_itm & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240
      & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_151_nl <= MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0(0)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(0)), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0(0)),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0(0)), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_0, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm(0)),
      STD_LOGIC_VECTOR'( and_1060_itm & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240
      & and_dcpl_207 & and_dcpl_847 & and_dcpl_583));
  not_5062_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_76_nl <= MUX1HOT_v_8_6_2((drf_output_sdt_2_sva_15_0_mx0w0(15
      DOWNTO 8)), attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_8, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_15_8,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_15_8, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_8, STD_LOGIC_VECTOR'(
      and_1062_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847));
  not_5088_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_136_nl <= MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0(7)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_7, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_7,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_7, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_7, STD_LOGIC_VECTOR'(
      and_1062_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_137_nl <= MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0(6)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_6, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_6,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_6, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_6, STD_LOGIC_VECTOR'(
      and_1062_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_138_nl <= MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0(5)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_5, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_5,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_5, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_5, STD_LOGIC_VECTOR'(
      and_1062_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_139_nl <= MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0(4)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_4, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_4,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_4, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_4, STD_LOGIC_VECTOR'(
      and_1062_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_140_nl <= MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0(3)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_3, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_3,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_3, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_3, STD_LOGIC_VECTOR'(
      and_1062_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_141_nl <= MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0(2)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_2, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_2,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_2, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_2, STD_LOGIC_VECTOR'(
      and_1062_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_142_nl <= MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0(1)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_1, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_1,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_1, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_1, STD_LOGIC_VECTOR'(
      and_1062_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847));
  attention_2_1_16_16_4_4_k_proj_re_mux1h_143_nl <= MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0(0)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_0, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_0,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_0, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_0, STD_LOGIC_VECTOR'(
      and_1062_ssc & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 &
      and_dcpl_847));
  and_1064_nl <= and_dcpl_732 AND and_dcpl_601;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_77_nl <= MUX1HOT_v_16_6_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_15_0, attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0, attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0_mx0w6,
      attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_15_0, STD_LOGIC_VECTOR'( and_1064_nl
      & and_dcpl_983 & and_dcpl_240 & and_dcpl_626 & and_dcpl_207 & and_dcpl_213));
  not_4571_nl <= NOT and_dcpl_619;
  nor_796_nl <= NOT((NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd) OR
      (NOT (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1))) OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2
      OR (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0)));
  mux_2038_nl <= MUX_s_1_2_2(mux_tmp_1945, mux_tmp_1943, nor_796_nl);
  and_1066_nl <= and_dcpl_732 AND and_dcpl_595;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_78_nl <= MUX1HOT_v_16_6_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_15_0,
      attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0, STD_LOGIC_VECTOR'( and_1066_nl
      & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847));
  not_4572_nl <= NOT and_dcpl_619;
  and_1420_nl <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1))
      AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 AND (NOT (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0)));
  mux_2039_nl <= MUX_s_1_2_2(mux_tmp_1945, mux_tmp_1943, and_1420_nl);
  and_1068_nl <= and_dcpl_732 AND and_dcpl_586;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_79_nl <= MUX1HOT_v_16_6_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_15_0,
      attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0, STD_LOGIC_VECTOR'( and_1068_nl
      & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847));
  not_4573_nl <= NOT and_dcpl_619;
  and_1613_nl <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1))
      AND (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2) AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0));
  mux_2040_nl <= MUX_s_1_2_2(mux_tmp_1945, mux_tmp_1943, and_1613_nl);
  and_1071_nl <= and_dcpl_732 AND and_dcpl_585 AND and_dcpl_462;
  and_1074_nl <= and_dcpl_743 AND and_dcpl_740 AND and_dcpl_854;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_80_nl <= MUX1HOT_v_16_8_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_15_0,
      attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0, output_0_15_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      STD_LOGIC_VECTOR'( and_1071_nl & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240
      & and_dcpl_207 & and_dcpl_847 & and_dcpl_739 & and_1074_nl));
  not_4574_nl <= NOT and_dcpl_619;
  or_2751_nl <= (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1))
      AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 AND (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0)))
      OR (NOT (fsm_output(6))) OR (fsm_output(8));
  and_1660_nl <= CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2=STD_LOGIC_VECTOR'("11"))
      AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd AND reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  mux_2045_nl <= MUX_s_1_2_2(mux_tmp_121, or_tmp_464, and_1660_nl);
  mux_2046_nl <= MUX_s_1_2_2(or_2751_nl, mux_2045_nl, fsm_output(4));
  mux_2047_nl <= MUX_s_1_2_2(or_tmp_464, mux_2046_nl, fsm_output(0));
  mux_2048_nl <= MUX_s_1_2_2(mux_2047_nl, mux_tmp_824, fsm_output(5));
  mux_2049_nl <= MUX_s_1_2_2(mux_2048_nl, mux_2025_cse, fsm_output(1));
  mux_2051_nl <= MUX_s_1_2_2(mux_2032_cse, mux_2049_nl, and_1773_cse);
  and_1075_nl <= and_dcpl_732 AND and_dcpl_598;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_81_nl <= MUX1HOT_v_16_6_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_15_0,
      attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0_mx0w1, STD_LOGIC_VECTOR'( and_1075_nl
      & attention_2_1_16_16_4_4_k_proj_re_or_cse & and_dcpl_983 & and_dcpl_240 &
      attention_2_1_16_16_4_4_k_proj_re_or_17_cse & and_dcpl_207));
  not_4575_nl <= NOT and_dcpl_619;
  or_2753_nl <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1/=STD_LOGIC_VECTOR'("01"))
      OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd;
  mux_2052_nl <= MUX_s_1_2_2(mux_tmp_1943, mux_tmp_1945, or_2753_nl);
  and_1081_nl <= and_dcpl_732 AND and_dcpl_610;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_82_nl <= MUX1HOT_v_16_6_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_15_0,
      attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0, STD_LOGIC_VECTOR'( and_1081_nl
      & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847));
  not_4576_nl <= NOT and_dcpl_619;
  or_2281_nl <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd OR (NOT (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1)))
      OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 OR (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0));
  mux_2053_nl <= MUX_s_1_2_2(mux_tmp_1943, mux_tmp_1945, or_2281_nl);
  and_1083_nl <= and_dcpl_732 AND and_dcpl_616;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_83_nl <= MUX1HOT_v_16_6_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_15_0,
      attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0, STD_LOGIC_VECTOR'( and_1083_nl
      & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847));
  not_4577_nl <= NOT and_dcpl_619;
  or_2292_nl <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd OR (NOT (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(1)))
      OR (NOT reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2) OR (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1(0));
  mux_2054_nl <= MUX_s_1_2_2(mux_tmp_1943, mux_tmp_1945, or_2292_nl);
  and_1086_nl <= and_dcpl_732 AND and_dcpl_591 AND and_dcpl_486;
  attention_2_1_16_16_4_4_k_proj_re_mux1h_84_nl <= MUX1HOT_v_16_6_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_15_0,
      attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0, STD_LOGIC_VECTOR'( and_1086_nl
      & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847));
  not_4578_nl <= NOT and_dcpl_619;
  or_2756_nl <= reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1/=STD_LOGIC_VECTOR'("11"))
      OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd;
  mux_2055_nl <= MUX_s_1_2_2(mux_tmp_1943, mux_tmp_1945, or_2756_nl);
  or_2757_nl <= CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("10"))
      OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  mux_2056_nl <= MUX_s_1_2_2(nor_1026_cse, mux_tmp_1578, or_2757_nl);
  and_1089_nl <= mux_2056_nl AND (NOT (fsm_output(8))) AND and_dcpl_814;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_51_nl <= MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_k_proj_re_0_2_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1,
      STD_LOGIC_VECTOR'( and_1089_nl & and_dcpl_989 & and_dcpl_374));
  not_4414_nl <= NOT and_dcpl_619;
  nor_1217_nl <= NOT((fsm_output(2)) OR reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      OR reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      OR reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 OR (NOT (fsm_output(4))));
  mux_2057_nl <= MUX_s_1_2_2(nor_1217_nl, and_1771_cse, fsm_output(1));
  and_1090_nl <= (fsm_output(0)) AND mux_2057_nl;
  mux_2058_nl <= MUX_s_1_2_2(and_1090_nl, (fsm_output(4)), fsm_output(3));
  or_3200_nl <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")) OR mux_2058_nl;
  or_3201_nl <= (NOT (fsm_output(6))) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_2059_nl <= MUX_s_1_2_2(or_3200_nl, or_3201_nl, fsm_output(5));
  attention_2_1_16_16_4_4_v_proj_re_mux1h_52_nl <= MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_k_proj_re_0_3_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1,
      STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16_mx0c1
      & and_dcpl_1003 & and_dcpl_207));
  not_4413_nl <= NOT and_dcpl_619;
  mux_2061_nl <= MUX_s_1_2_2(and_dcpl_364, and_1771_cse, fsm_output(1));
  or_2763_nl <= (fsm_output(5)) OR ((fsm_output(0)) AND mux_2061_nl);
  mux_2062_nl <= MUX_s_1_2_2(or_2763_nl, or_2699_cse, fsm_output(3));
  or_2764_nl <= (fsm_output(6)) OR mux_2062_nl;
  mux_2063_nl <= MUX_s_1_2_2(not_tmp_253, or_2764_nl, fsm_output(7));
  or_2765_nl <= reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 OR CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd/=STD_LOGIC_VECTOR'("001"));
  mux_2064_nl <= MUX_s_1_2_2(or_1983_cse, mux_tmp_1562, or_2765_nl);
  and_1097_nl <= (NOT(mux_2064_nl OR (fsm_output(8)))) AND and_dcpl_748;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_53_nl <= MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_q_proj_re_0_2_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1,
      STD_LOGIC_VECTOR'( and_1097_nl & and_dcpl_999 & and_dcpl_374));
  not_4412_nl <= NOT and_dcpl_619;
  nand_370_nl <= NOT((NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))))
      AND (fsm_output(4)));
  mux_2065_nl <= MUX_s_1_2_2(nand_370_nl, or_tmp_330, fsm_output(3));
  mux_2068_nl <= MUX_s_1_2_2(mux_tmp_2067, mux_2065_nl, or_1880_cse);
  attention_2_1_16_16_4_4_v_proj_re_mux1h_54_nl <= MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_q_proj_re_0_3_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg(39 DOWNTO 16)), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1,
      STD_LOGIC_VECTOR'( apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16_mx0c1
      & and_dcpl_959 & and_dcpl_207));
  not_nl <= NOT and_dcpl_619;
  attention_2_1_16_16_4_4_v_proj_re_mux1h_55_nl <= MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_v_proj_re_0_4_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_39_16, RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      STD_LOGIC_VECTOR'( and_dcpl_726 & and_dcpl_410 & and_dcpl_240));
  not_4579_nl <= NOT and_dcpl_619;
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_36_nl <= MUX_v_24_16_2(attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_39_16, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  attention_2_1_16_16_4_4_v_proj_re_mux1h_56_nl <= MUX1HOT_v_24_9_2(attention_2_1_16_16_4_4_v_proj_re_0_13_sva_1_39_16,
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48_mx0w2, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_39_16, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16_mx0w1,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16_mx0w1,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_36_nl, LINEAR_FORWARD_NO_MUL_LOOP_2_3_conc_1_mut_71_48_mx0w3,
      STD_LOGIC_VECTOR'( and_dcpl_726 & and_dcpl_257 & attention_2_1_16_16_4_4_k_proj_re_or_cse
      & and_dcpl_983 & and_dcpl_240 & attention_2_1_16_16_4_4_k_proj_re_or_17_cse
      & and_dcpl_207 & and_dcpl_583 & and_dcpl_265));
  not_4580_nl <= NOT and_dcpl_619;
  LINEAR_FORWARD_NO_MUL_LOOP_2_mux_33_nl <= MUX_v_24_16_2(attention_2_1_16_16_4_4_q_proj_re_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_1_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_re_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_3_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_re_0_4_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_5_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_re_0_6_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_7_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_re_0_8_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_9_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_re_0_10_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_11_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_re_0_12_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_13_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_re_0_14_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_15_sva_1_39_16, reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
      & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_38_nl <= MUX_v_24_16_2(attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_39_16,
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  attention_2_1_16_16_4_4_v_proj_re_mux1h_57_nl <= MUX1HOT_v_24_8_2(attention_2_1_16_16_4_4_v_proj_re_0_11_sva_1_39_16,
      LINEAR_FORWARD_NO_MUL_LOOP_2_mux_33_nl, attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_39_16, attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16_mx0w1,
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16_mx0w1, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_38_nl, STD_LOGIC_VECTOR'( and_dcpl_726 & and_dcpl_257
      & and_dcpl_1011 & and_dcpl_983 & and_dcpl_240 & and_dcpl_207 & and_dcpl_847
      & and_dcpl_583));
  not_4581_nl <= NOT and_dcpl_619;
  QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_nl
      <= NOT((NOT QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1)
      OR QUANTIZE_ACTIVATION_LOOP_3_nand_seb);
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_nl <= MUX_v_8_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(15
      DOWNTO 8)), (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1(15 DOWNTO
      8)), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_15_8, apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_8,
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3(15 DOWNTO 8)), (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm(15
      DOWNTO 8)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_8, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3(15
      DOWNTO 8)), (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm(15 DOWNTO
      8)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_13
      & apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_12_8), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3(15
      DOWNTO 8)), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm(15 DOWNTO
      8)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_8,
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_nl <= MUX_v_8_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(15
      DOWNTO 8)), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_8, attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_8,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_ftd, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_15_8,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(15 DOWNTO 8)), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_13
      & (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(12 DOWNTO 8))), attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_8,
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(15 DOWNTO 8)), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(15
      DOWNTO 8)), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0(15 DOWNTO 8)),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0(15 DOWNTO 8)), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(15
      DOWNTO 8)), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(15 DOWNTO 8)),
      (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0(15 DOWNTO 8)), (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0(15
      DOWNTO 8)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_66_nl <= MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(7)),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1(7)), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_7,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_7, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3(7)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm(7)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_7, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3(7)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm(7)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_7, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3(7)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm(7)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_7, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_74_nl <= MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(6)),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1(6)), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_6,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_6, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3(6)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm(6)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_2,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_6, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3(6)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm(6)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_2,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_6, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3(6)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm(6)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_2,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_6, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_75_nl <= MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(5)),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1(5)), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_5,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_5, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3(5)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm(5)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_3,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_5, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3(5)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm(5)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_3,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_5, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3(5)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm(5)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_3,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_5, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_76_nl <= MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(4)),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1(4)), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_4,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_4, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3(4)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm(4)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_4,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_4, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3(4)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm(4)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_4,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_4, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3(4)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm(4)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_4,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_4, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_77_nl <= MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(3)),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1(3)), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_3,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_3, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3(3)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm(3)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_5,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_3, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3(3)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm(3)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_5,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_3, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3(3)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm(3)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_5,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_3, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_78_nl <= MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(2)),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1(2)), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_2,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_2, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3(2)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm(2)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_6,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_2, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3(2)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm(2)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_6,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_2, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3(2)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm(2)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_6,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_2, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_79_nl <= MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(1)),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1(1)), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_1, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3(1)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm(1)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_7,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_1, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3(1)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm(1)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_7,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_1, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3(1)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm(1)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_7,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_1, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_80_nl <= MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(0)),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1(0)), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_0,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_0, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3(0)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm(0)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_8,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_0, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3(0)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm(0)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_8,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_0, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3(0)),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm(0)), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_8,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_0, STD_LOGIC_VECTOR'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_61_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(7)),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_7, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_7,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(7)), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(7)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_7, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(7)),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(7)), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0(7)),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0(7)), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(7)),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(7)), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0(7)),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0(7)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_81_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(6)),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_6, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_1,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_1, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_6,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(6)), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(6)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_6, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(6)),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(6)), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0(6)),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0(6)), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(6)),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(6)), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0(6)),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0(6)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_82_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(5)),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_5, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_2,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_2, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_5,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(5)), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(5)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_5, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(5)),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(5)), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0(5)),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0(5)), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(5)),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(5)), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0(5)),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0(5)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_83_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(4)),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_4, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_3,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_3, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_4,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(4)), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(4)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_4, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(4)),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(4)), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0(4)),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0(4)), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(4)),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(4)), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0(4)),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0(4)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_84_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(3)),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_3, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_4,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_4, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_3,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(3)), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(3)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_3, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(3)),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(3)), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0(3)),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0(3)), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(3)),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(3)), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0(3)),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0(3)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_85_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(2)),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_2, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_5,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_5, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_2,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(2)), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(2)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_2, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(2)),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(2)), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0(2)),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0(2)), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(2)),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(2)), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0(2)),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0(2)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_86_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(1)),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_1, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_6,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_6, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_1,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(1)), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(1)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_1, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(1)),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(1)), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0(1)),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0(1)), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(1)),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(1)), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0(1)),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0(1)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_87_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0(0)),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_0, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_7,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_7, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_0,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0(0)), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0(0)),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_0, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0(0)),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0(0)), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0(0)),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0(0)), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0(0)),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0(0)), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0(0)),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0(0)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_32_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(15)),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(15)), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(15)),
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_15, (attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8(7)),
      (attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8(7)), (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8(7)),
      (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8(7)), (attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8(7)),
      (attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8(7)), (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8(7)),
      (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8(7)), (attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8(7)),
      (attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8(7)), (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8(7)),
      (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8(7)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_70_nl <= MUX_v_3_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(14
      DOWNTO 12)), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(14 DOWNTO 12)),
      (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(14 DOWNTO 12)), attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_14_12,
      (attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8(6 DOWNTO 4)), (attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8(6
      DOWNTO 4)), (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8(6 DOWNTO 4)),
      (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8(6 DOWNTO 4)), (attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8(6
      DOWNTO 4)), (attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8(6 DOWNTO 4)),
      (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8(6 DOWNTO 4)), (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8(6
      DOWNTO 4)), (attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8(6 DOWNTO 4)),
      (attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8(6 DOWNTO 4)), (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8(6
      DOWNTO 4)), (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8(6 DOWNTO 4)),
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_71_nl <= MUX_v_3_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(11
      DOWNTO 9)), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(11 DOWNTO 9)),
      (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(11 DOWNTO 9)), attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_11_9,
      (attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8(3 DOWNTO 1)), (attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8(3
      DOWNTO 1)), (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8(3 DOWNTO 1)),
      (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8(3 DOWNTO 1)), (attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8(3
      DOWNTO 1)), (attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8(3 DOWNTO 1)),
      (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8(3 DOWNTO 1)), (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8(3
      DOWNTO 1)), (attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8(3 DOWNTO 1)),
      (attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8(3 DOWNTO 1)), (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8(3
      DOWNTO 1)), (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8(3 DOWNTO 1)),
      STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_72_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(8)),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(8)), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(8)),
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_8, (attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8(0)),
      (attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8(0)), (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8(0)),
      (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8(0)), (attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8(0)),
      (attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8(0)), (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8(0)),
      (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8(0)), (attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8(0)),
      (attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8(0)), (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8(0)),
      (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8(0)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_50_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(7)),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(7)), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(7)),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(7)), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_7, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_7, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_7, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_7, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_7, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_7, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_51_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(6)),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(6)), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(6)),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(6)), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_6, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_6, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_6, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_6, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_6, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_6, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_52_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(5)),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(5)), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(5)),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(5)), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_5, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_5, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_5, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_5, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_5, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_5, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_53_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(4)),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(4)), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(4)),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(4)), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_4, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_4, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_4, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_4, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_4, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_4, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_54_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(3)),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(3)), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(3)),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(3)), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_3, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_3, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_3, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_3, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_3, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_3, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_55_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(2)),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(2)), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(2)),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(2)), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_2, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_2, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_2, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_2, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_2, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_2, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_56_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(1)),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(1)), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(1)),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(1)), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_1, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_1, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_1, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_1, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_1, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_1, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux_57_nl <= MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0(0)),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0(0)), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0(0)),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0(0)), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_0, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_0, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_0, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_0, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_0, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_0, STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1));
  APPLY_ROTARY_POS_EMB_LOOP_3_and_7_nl <= (NOT reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1)
      AND reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  APPLY_ROTARY_POS_EMB_LOOP_3_and_5_nl <= reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      AND reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  mux_2129_nl <= MUX_s_1_2_2((NOT and_1570_cse), or_tmp_762, fsm_output(5));
  mux_2130_nl <= MUX_s_1_2_2(mux_2129_nl, or_tmp_682, fsm_output(3));
  mux_2131_nl <= MUX_s_1_2_2(and_1559_cse, (NOT or_3137_cse), fsm_output(3));
  attention_2_1_16_16_4_4_q_embed_or_nl <= attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c1
      OR (or_dcpl_996 AND and_dcpl_204);
  attention_2_1_16_16_4_4_q_embed_and_33_nl <= (NOT or_dcpl_996) AND and_dcpl_204;
  attention_2_1_16_16_4_4_q_embed_mux1h_40_nl <= MUX1HOT_v_40_9_2(attention_2_1_16_16_4_4_q_embed_0_0_2_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1, APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2, attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx1,
      attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx2, attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1,
      (ATTN_2D_LOOP_3_mux_16_itm & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( and_dcpl_346 & attention_2_1_16_16_4_4_q_embed_or_nl & attention_2_1_16_16_4_4_q_embed_and_33_nl
      & and_dcpl_348 & and_dcpl_349 & and_dcpl_351 & and_dcpl_1162 & and_dcpl_352
      & attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c9));
  not_4510_nl <= NOT mux_tmp_2153;
  attention_2_1_16_16_4_4_q_embed_mux1h_41_nl <= MUX1HOT_v_40_6_2(attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1,
      attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2,
      attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx1, (ATTN_2D_LOOP_3_mux_16_itm
      & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( and_dcpl_346 & and_dcpl_204 & and_dcpl_348 & and_dcpl_351
      & and_dcpl_352 & attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx0c7));
  not_4483_nl <= NOT mux_tmp_2176;
  nor_1245_nl <= NOT((NOT(CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)/=STD_LOGIC_VECTOR'("00")) OR reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 OR
      (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0))) OR CONV_SL_1_1(fsm_output(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10111")))) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_2158_nl <= MUX_s_1_2_2(mux_2157_cse, nor_1245_nl, fsm_output(5));
  mux_2159_nl <= MUX_s_1_2_2(nor_1239_cse, mux_2158_nl, fsm_output(7));
  attention_2_1_16_16_4_4_q_embed_mux1h_42_nl <= MUX1HOT_v_40_6_2(attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1,
      attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2,
      attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx1, (ATTN_2D_LOOP_3_mux_16_itm
      & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( and_dcpl_346 & and_dcpl_204 & and_dcpl_348 & and_dcpl_351
      & and_dcpl_352 & attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx0c7));
  not_4482_nl <= NOT mux_tmp_2176;
  nor_1256_nl <= NOT((NOT(CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)/=STD_LOGIC_VECTOR'("00")) OR (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1)
      OR (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0))) OR CONV_SL_1_1(fsm_output(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10111")))) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_2181_nl <= MUX_s_1_2_2(mux_2157_cse, nor_1256_nl, fsm_output(5));
  mux_2182_nl <= MUX_s_1_2_2(nor_1239_cse, mux_2181_nl, fsm_output(7));
  attention_2_1_16_16_4_4_q_embed_or_5_nl <= attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c1
      OR (or_dcpl_988 AND and_dcpl_204);
  attention_2_1_16_16_4_4_q_embed_and_35_nl <= (NOT or_dcpl_988) AND and_dcpl_204;
  attention_2_1_16_16_4_4_q_embed_mux1h_43_nl <= MUX1HOT_v_40_9_2(attention_2_1_16_16_4_4_q_embed_1_0_1_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1, APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2, attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx1,
      attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx2, attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1,
      (ATTN_2D_LOOP_3_mux_16_itm & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( and_dcpl_346 & attention_2_1_16_16_4_4_q_embed_or_5_nl &
      attention_2_1_16_16_4_4_q_embed_and_35_nl & and_dcpl_348 & and_dcpl_349 & and_dcpl_351
      & and_dcpl_1162 & and_dcpl_352 & attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c9));
  not_4511_nl <= NOT mux_tmp_2153;
  attention_2_1_16_16_4_4_q_embed_mux1h_44_nl <= MUX1HOT_v_40_6_2(attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1,
      attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2,
      attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx1, (ATTN_2D_LOOP_3_mux_16_itm
      & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( and_dcpl_346 & and_dcpl_204 & and_dcpl_348 & and_dcpl_351
      & and_dcpl_352 & attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx0c7));
  not_4512_nl <= NOT mux_tmp_2176;
  nor_1272_nl <= NOT((NOT(CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)/=STD_LOGIC_VECTOR'("01")) OR (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1)
      OR (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0)) OR CONV_SL_1_1(fsm_output(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10111")))) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_2197_nl <= MUX_s_1_2_2(mux_2157_cse, nor_1272_nl, fsm_output(5));
  mux_2198_nl <= MUX_s_1_2_2(nor_1239_cse, mux_2197_nl, fsm_output(7));
  attention_2_1_16_16_4_4_q_embed_mux1h_45_nl <= MUX1HOT_v_40_6_2(attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1,
      attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2,
      attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx1, (ATTN_2D_LOOP_3_mux_16_itm
      & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( and_dcpl_346 & and_dcpl_204 & and_dcpl_348 & and_dcpl_351
      & and_dcpl_352 & attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx0c7));
  not_4513_nl <= NOT mux_tmp_2176;
  nor_1283_nl <= NOT((NOT(CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)/=STD_LOGIC_VECTOR'("01")) OR reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 OR
      (NOT (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0))) OR CONV_SL_1_1(fsm_output(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10111")))) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_2203_nl <= MUX_s_1_2_2(mux_2157_cse, nor_1283_nl, fsm_output(5));
  mux_2204_nl <= MUX_s_1_2_2(nor_1239_cse, mux_2203_nl, fsm_output(7));
  attention_2_1_16_16_4_4_q_embed_mux1h_46_nl <= MUX1HOT_v_40_6_2(attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1,
      attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2,
      attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx1, (ATTN_2D_LOOP_3_mux_16_itm
      & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( and_dcpl_346 & and_dcpl_204 & and_dcpl_348 & and_dcpl_351
      & and_dcpl_352 & attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx0c7));
  not_4514_nl <= NOT mux_tmp_2176;
  nor_1294_nl <= NOT((CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)=STD_LOGIC_VECTOR'("01")) AND reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 AND
      (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0)) AND CONV_SL_1_1(fsm_output(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("10111"))) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_2209_nl <= MUX_s_1_2_2(mux_2157_cse, nor_1294_nl, fsm_output(5));
  mux_2210_nl <= MUX_s_1_2_2(nor_1239_cse, mux_2209_nl, fsm_output(7));
  attention_2_1_16_16_4_4_q_embed_or_6_nl <= attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c1
      OR (or_dcpl_987 AND and_dcpl_204);
  attention_2_1_16_16_4_4_q_embed_and_37_nl <= (NOT or_dcpl_987) AND and_dcpl_204;
  attention_2_1_16_16_4_4_q_embed_mux1h_47_nl <= MUX1HOT_v_40_9_2(attention_2_1_16_16_4_4_q_embed_2_0_1_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1, APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2, attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx1,
      attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx2, attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1,
      (ATTN_2D_LOOP_3_mux_16_itm & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( and_dcpl_346 & attention_2_1_16_16_4_4_q_embed_or_6_nl &
      attention_2_1_16_16_4_4_q_embed_and_37_nl & and_dcpl_348 & and_dcpl_349 & and_dcpl_351
      & and_dcpl_1162 & and_dcpl_352 & attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c9));
  not_4515_nl <= NOT mux_tmp_2153;
  attention_2_1_16_16_4_4_q_embed_mux1h_48_nl <= MUX1HOT_v_40_6_2(attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1,
      attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2,
      attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx1, (ATTN_2D_LOOP_3_mux_16_itm
      & ATTN_2D_LOOP_3_mux_17_itm), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      STD_LOGIC_VECTOR'( and_dcpl_346 & and_dcpl_204 & and_dcpl_348 & and_dcpl_351
      & and_dcpl_352 & attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx0c7));
  not_4516_nl <= NOT mux_tmp_2176;
  nor_1310_nl <= NOT((NOT(CONV_SL_1_1(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2 DOWNTO
      1)/=STD_LOGIC_VECTOR'("10")) OR (NOT reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1)
      OR (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0)) OR CONV_SL_1_1(fsm_output(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10111")))) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_2225_nl <= MUX_s_1_2_2(mux_2157_cse, nor_1310_nl, fsm_output(5));
  mux_2226_nl <= MUX_s_1_2_2(nor_1239_cse, mux_2225_nl, fsm_output(7));
  GEMM_3D_FLOAT_LOOP_3_not_28_nl <= NOT GEMM_3D_FLOAT_LOOP_3_and_tmp_sva_mx0w0;
  GEMM_3D_FLOAT_LOOP_3_and_35_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1, GEMM_3D_FLOAT_LOOP_3_not_28_nl);
  GEMM_3D_FLOAT_LOOP_3_not_27_nl <= NOT GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva_mx0w0;
  GEMM_3D_FLOAT_LOOP_3_and_34_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1, GEMM_3D_FLOAT_LOOP_3_not_27_nl);
  GEMM_3D_FLOAT_LOOP_3_not_26_nl <= NOT GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva_mx0w0;
  GEMM_3D_FLOAT_LOOP_3_and_33_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1, GEMM_3D_FLOAT_LOOP_3_not_26_nl);
  GEMM_3D_FLOAT_LOOP_3_not_25_nl <= NOT GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva_mx0w0;
  GEMM_3D_FLOAT_LOOP_3_and_32_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1, GEMM_3D_FLOAT_LOOP_3_not_25_nl);
  GEMM_3D_FLOAT_LOOP_3_not_24_nl <= NOT GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva_mx0w0;
  GEMM_3D_FLOAT_LOOP_3_and_31_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1, GEMM_3D_FLOAT_LOOP_3_not_24_nl);
  GEMM_3D_FLOAT_LOOP_3_not_23_nl <= NOT GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva_mx0w0;
  GEMM_3D_FLOAT_LOOP_3_and_30_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1, GEMM_3D_FLOAT_LOOP_3_not_23_nl);
  GEMM_3D_FLOAT_LOOP_3_not_22_nl <= NOT GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva_mx0w0;
  GEMM_3D_FLOAT_LOOP_3_and_29_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1, GEMM_3D_FLOAT_LOOP_3_not_22_nl);
  GEMM_3D_FLOAT_LOOP_3_not_21_nl <= NOT GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva_mx0w0;
  GEMM_3D_FLOAT_LOOP_3_and_28_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1, GEMM_3D_FLOAT_LOOP_3_not_21_nl);
  GEMM_3D_FLOAT_LOOP_3_not_20_nl <= NOT GEMM_3D_FLOAT_LOOP_3_and_tmp_4_sva_mx0w2;
  GEMM_3D_FLOAT_LOOP_3_and_27_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1, GEMM_3D_FLOAT_LOOP_3_not_20_nl);
  GEMM_3D_FLOAT_LOOP_3_not_19_nl <= NOT GEMM_3D_FLOAT_LOOP_3_and_tmp_7_sva_mx0w1;
  GEMM_3D_FLOAT_LOOP_3_and_26_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1, GEMM_3D_FLOAT_LOOP_3_not_19_nl);
  GEMM_3D_FLOAT_LOOP_3_not_18_nl <= NOT GEMM_3D_FLOAT_LOOP_3_and_tmp_5_sva_mx0w2;
  GEMM_3D_FLOAT_LOOP_3_and_25_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1, GEMM_3D_FLOAT_LOOP_3_not_18_nl);
  GEMM_3D_FLOAT_LOOP_3_not_17_nl <= NOT GEMM_3D_FLOAT_LOOP_3_and_tmp_6_sva_mx0w1;
  GEMM_3D_FLOAT_LOOP_3_and_24_nl <= MUX_v_40_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000"),
      attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1, GEMM_3D_FLOAT_LOOP_3_not_17_nl);
  nor_1319_nl <= NOT((fsm_output(3)) OR (fsm_output(5)) OR or_tmp_1632);
  mux_2248_nl <= MUX_s_1_2_2(mux_tmp_857, nor_1319_nl, fsm_output(6));
  output_and_35_nl <= or_dcpl_1155 AND (NOT and_dcpl_1232);
  output_and_39_nl <= or_dcpl_1158 AND (NOT and_dcpl_1232);
  output_and_43_nl <= or_dcpl_1160 AND (NOT and_dcpl_1232);
  output_and_47_nl <= or_dcpl_1162 AND (NOT and_dcpl_1232);
  output_and_51_nl <= or_dcpl_1165 AND (NOT and_dcpl_1232);
  output_and_55_nl <= or_dcpl_1167 AND (NOT and_dcpl_1232);
  output_and_59_nl <= or_dcpl_1169 AND (NOT and_dcpl_1232);
  output_and_63_nl <= or_dcpl_1141 AND (NOT and_dcpl_1232);
  output_and_61_nl <= or_dcpl_1170 AND (NOT and_dcpl_1232);
  output_and_57_nl <= or_dcpl_1168 AND (NOT and_dcpl_1232);
  output_and_53_nl <= or_dcpl_1166 AND (NOT and_dcpl_1232);
  output_and_49_nl <= or_dcpl_1164 AND (NOT and_dcpl_1232);
  output_and_45_nl <= or_dcpl_1161 AND (NOT and_dcpl_1232);
  output_and_41_nl <= or_dcpl_1159 AND (NOT and_dcpl_1232);
  output_and_37_nl <= or_dcpl_1156 AND (NOT and_dcpl_1232);
  output_and_33_nl <= or_dcpl_1152 AND (NOT and_dcpl_1232);
  GEMM_3D_FLOAT_LOOP_4_l_mux1h_6_nl <= MUX1HOT_s_1_3_2((z_out_3(1)), (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_k_2_0_sva_1(1)),
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(1)), STD_LOGIC_VECTOR'(
      GEMM_3D_FLOAT_LOOP_4_l_or_2_cse & GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c3
      & and_dcpl_193));
  operator_40_24_true_AC_TRN_AC_WRAP_or_nl <= CONV_SL_1_1(acc_3_cse_40_1(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0000"));
  compute_sqrt_for_acc_3_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(z_out_12(3
      DOWNTO 1)), 3), 4) + SIGNED'( "1011"), 4));
  RMS_NORM_LOOP_2_and_35_nl <= RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_mux1h_itm AND (NOT(RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_nor_1_ssc_1
      OR RMS_NORM_LOOP_2_and_33_ssc_1));
  nor_658_nl <= NOT(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 OR reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1);
  RMS_NORM_LOOP_2_2_and_35_nl <= RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_mux1h_itm AND
      (NOT(RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_nor_1_ssc_1 OR RMS_NORM_LOOP_2_2_and_33_ssc_1));
  mux_1258_nl <= MUX_s_1_2_2(or_tmp_1664, mux_tmp_1245, and_1559_cse);
  mux_1254_nl <= MUX_s_1_2_2(or_tmp_1066, mux_tmp_1237, fsm_output(5));
  mux_1255_nl <= MUX_s_1_2_2(mux_1254_nl, mux_tmp_1250, fsm_output(0));
  mux_1256_nl <= MUX_s_1_2_2(mux_tmp_1245, mux_1255_nl, fsm_output(2));
  or_2167_nl <= (fsm_output(8)) OR mux_792_cse;
  mux_1252_nl <= MUX_s_1_2_2(or_2167_nl, or_1197_cse, fsm_output(5));
  mux_1247_nl <= MUX_s_1_2_2(or_tmp_1066, or_1984_cse, fsm_output(5));
  mux_1251_nl <= MUX_s_1_2_2(mux_tmp_1250, mux_1247_nl, fsm_output(0));
  mux_1253_nl <= MUX_s_1_2_2(mux_1252_nl, mux_1251_nl, fsm_output(2));
  mux_1257_nl <= MUX_s_1_2_2(mux_1256_nl, mux_1253_nl, fsm_output(1));
  mux_1259_nl <= MUX_s_1_2_2(mux_1258_nl, mux_1257_nl, fsm_output(4));
  or_3075_nl <= (fsm_output(0)) OR (fsm_output(2));
  mux_1243_nl <= MUX_s_1_2_2(mux_tmp_1240, mux_tmp_1238, or_3075_nl);
  nor_374_nl <= NOT(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd OR reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      OR CONV_SL_1_1(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(0))));
  mux_1241_nl <= MUX_s_1_2_2(mux_tmp_1238, mux_tmp_1240, nor_374_nl);
  or_2162_nl <= (fsm_output(5)) OR mux_tmp_1237;
  mux_1239_nl <= MUX_s_1_2_2(mux_tmp_1238, or_2162_nl, fsm_output(0));
  mux_1242_nl <= MUX_s_1_2_2(mux_1241_nl, mux_1239_nl, fsm_output(2));
  mux_1244_nl <= MUX_s_1_2_2(mux_1243_nl, mux_1242_nl, fsm_output(1));
  mux_1246_nl <= MUX_s_1_2_2(mux_tmp_1245, mux_1244_nl, fsm_output(4));
  mux_1260_nl <= MUX_s_1_2_2(mux_1259_nl, mux_1246_nl, fsm_output(3));
  operator_40_24_true_AC_TRN_AC_WRAP_mux1h_nl <= MUX1HOT_s_1_7_2(operator_40_24_true_AC_TRN_AC_WRAP_or_nl,
      (compute_sqrt_for_acc_3_nl(3)), reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1,
      RMS_NORM_LOOP_2_and_35_nl, nor_658_nl, RMS_NORM_LOOP_2_2_and_35_nl, (NOT QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1),
      STD_LOGIC_VECTOR'( rms_norm_16_variance_or_1_cse & and_dcpl_382 & (NOT mux_1260_nl)
      & and_dcpl_344 & and_dcpl_207 & and_dcpl_548 & and_dcpl_557));
  nor_1048_nl <= NOT((fsm_output(5)) OR (fsm_output(0)) OR (NOT (fsm_output(4))));
  and_1603_nl <= (fsm_output(5)) AND (fsm_output(0)) AND (fsm_output(1)) AND (NOT
      (fsm_output(4)));
  mux_1261_nl <= MUX_s_1_2_2(nor_1048_nl, and_1603_nl, fsm_output(3));
  QUANTIZE_ACTIVATION_LOOP_1_1_max_val_asn_GEMM_3D_FLOAT_LOOP_4_l_2_operator_40_24_true_AC_TRN_AC_WRAP_or_nl
      <= (operator_40_24_true_AC_TRN_AC_WRAP_mux1h_nl AND (NOT(mux_1261_nl AND and_dcpl_390)))
      OR and_dcpl_442;
  and_1256_nl <= and_dcpl_191 AND mux_tmp_787 AND and_dcpl_293;
  mux_2246_nl <= MUX_s_1_2_2(and_1762_cse, and_tmp_42, fsm_output(3));
  nor_1318_nl <= NOT((fsm_output(3)) OR (fsm_output(5)) OR mux_tmp_1281);
  mux_2247_nl <= MUX_s_1_2_2(mux_2246_nl, nor_1318_nl, fsm_output(6));
  and_1257_nl <= mux_2247_nl AND GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c6;
  GEMM_3D_FLOAT_LOOP_4_l_mux1h_8_nl <= MUX1HOT_s_1_7_2(QUANTIZE_ACTIVATION_LOOP_1_1_max_val_asn_GEMM_3D_FLOAT_LOOP_4_l_2_operator_40_24_true_AC_TRN_AC_WRAP_or_nl,
      (z_out_3(0)), (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_k_2_0_sva_1(0)), (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0)),
      CACHE_UPDATE_LOOP_2_1_acc_2_itm_2_1, reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1,
      CACHE_UPDATE_LOOP_2_acc_2_itm_2_1, STD_LOGIC_VECTOR'( GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c0
      & GEMM_3D_FLOAT_LOOP_4_l_or_2_cse & GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c3
      & and_dcpl_193 & and_1256_nl & and_1257_nl & and_dcpl_316));
  CACHE_UPDATE_LOOP_3_mux1h_6_nl <= MUX1HOT_s_1_3_2(reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0,
      reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd, (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(1)),
      STD_LOGIC_VECTOR'( CACHE_UPDATE_LOOP_3_or_cse & CACHE_UPDATE_LOOP_3_or_1_cse
      & and_dcpl_1294));
  CACHE_UPDATE_LOOP_3_mux1h_7_nl <= MUX1HOT_s_1_3_2(reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1,
      reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1, (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0)),
      STD_LOGIC_VECTOR'( CACHE_UPDATE_LOOP_3_or_cse & CACHE_UPDATE_LOOP_3_or_1_cse
      & and_dcpl_1294));
  z_out_3 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'(
      CACHE_UPDATE_LOOP_3_mux1h_6_nl & CACHE_UPDATE_LOOP_3_mux1h_7_nl), 2), 3) +
      UNSIGNED'( "001"), 3));
  z_out_4 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'(
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1),
      2), 3) + UNSIGNED'( "001"), 3));
  GEMM_3D_FLOAT_LOOP_1_GEMM_3D_FLOAT_LOOP_1_mux_2_nl <= MUX_s_1_2_2(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd, GEMM_3D_FLOAT_LOOP_1_or_ssc);
  GEMM_3D_FLOAT_LOOP_1_GEMM_3D_FLOAT_LOOP_1_mux_3_nl <= MUX_s_1_2_2(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1, GEMM_3D_FLOAT_LOOP_1_or_ssc);
  z_out_5 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'(
      GEMM_3D_FLOAT_LOOP_1_GEMM_3D_FLOAT_LOOP_1_mux_2_nl & GEMM_3D_FLOAT_LOOP_1_GEMM_3D_FLOAT_LOOP_1_mux_3_nl),
      2), 3) + UNSIGNED'( "001"), 3));
  acc_3_cse_40_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1) + UNSIGNED(reg_RMS_NORM_LOOP_1_1_slc_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_mul_55_16_cse_1_slc
      & (APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm(39 DOWNTO 16))), 40));
  APPLY_ROTARY_POS_EMB_LOOP_6_APPLY_ROTARY_POS_EMB_LOOP_6_or_8_nl <= (NOT(and_dcpl_1371
      OR and_dcpl_1379)) OR and_dcpl_1385;
  APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_36_nl <= MUX1HOT_v_13_3_2(reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1,
      STD_LOGIC_VECTOR'( "0110100011101"), STD_LOGIC_VECTOR'( "1110001000111"), STD_LOGIC_VECTOR'(
      and_dcpl_1371 & and_dcpl_1379 & and_dcpl_1385));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_37_nl <= MUX1HOT_v_24_3_2(for_for_strm_in_tmp_sva_25_2,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(39 DOWNTO 16)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(39
      DOWNTO 16)), STD_LOGIC_VECTOR'( and_dcpl_1371 & and_dcpl_1379 & and_dcpl_1385));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_38_nl <= MUX1HOT_v_8_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(15 DOWNTO 8)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(15
      DOWNTO 8)), STD_LOGIC_VECTOR'( and_dcpl_1371 & and_dcpl_1379 & and_dcpl_1385));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_39_nl <= MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(7)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(7)),
      STD_LOGIC_VECTOR'( and_dcpl_1371 & and_dcpl_1379 & and_dcpl_1385));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_40_nl <= MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(6)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(6)),
      STD_LOGIC_VECTOR'( and_dcpl_1371 & and_dcpl_1379 & and_dcpl_1385));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_41_nl <= MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(5)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(5)),
      STD_LOGIC_VECTOR'( and_dcpl_1371 & and_dcpl_1379 & and_dcpl_1385));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_42_nl <= MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(4)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(4)),
      STD_LOGIC_VECTOR'( and_dcpl_1371 & and_dcpl_1379 & and_dcpl_1385));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_43_nl <= MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(3)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(3)),
      STD_LOGIC_VECTOR'( and_dcpl_1371 & and_dcpl_1379 & and_dcpl_1385));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_44_nl <= MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(2)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(2)),
      STD_LOGIC_VECTOR'( and_dcpl_1371 & and_dcpl_1379 & and_dcpl_1385));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_45_nl <= MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(1)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(1)),
      STD_LOGIC_VECTOR'( and_dcpl_1371 & and_dcpl_1379 & and_dcpl_1385));
  APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_46_nl <= MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(0)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(0)),
      STD_LOGIC_VECTOR'( and_dcpl_1371 & and_dcpl_1379 & and_dcpl_1385));
  z_out_9 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( CONV_SIGNED(CONV_UNSIGNED(UNSIGNED((NOT
      and_dcpl_1371) & '0' & (NOT and_dcpl_1371) & APPLY_ROTARY_POS_EMB_LOOP_6_APPLY_ROTARY_POS_EMB_LOOP_6_or_8_nl
      & (NOT and_dcpl_1385) & (NOT and_dcpl_1385) & (NOT and_dcpl_1385) & APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_36_nl),
      20), 21) * SIGNED(APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_37_nl & APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_38_nl
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_39_nl & APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_40_nl
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_41_nl & APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_42_nl
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_43_nl & APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_44_nl
      & APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_45_nl & APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_46_nl)),
      60));
  RMS_NORM_LOOP_1_1_mux1h_134_nl <= MUX1HOT_s_1_4_2((for_for_strm_in_tmp_sva_31_26(5)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(39)), QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39,
      (APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16(23)), STD_LOGIC_VECTOR'( and_dcpl_1393
      & RMS_NORM_LOOP_1_1_or_3_ssc & RMS_NORM_LOOP_1_1_or_1_ssc & and_dcpl_1415));
  RMS_NORM_LOOP_1_1_and_14_nl <= RMS_NORM_LOOP_1_1_mux1h_134_nl AND RMS_NORM_LOOP_1_1_nor_seb;
  RMS_NORM_LOOP_1_1_mux1h_135_nl <= MUX1HOT_v_3_4_2(STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(for_for_strm_in_tmp_sva_31_26(5),
      1),3)), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(38 DOWNTO 36)), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(38
      DOWNTO 36)), (APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16(22 DOWNTO 20)),
      STD_LOGIC_VECTOR'( and_dcpl_1393 & RMS_NORM_LOOP_1_1_or_3_ssc & RMS_NORM_LOOP_1_1_or_1_ssc
      & and_dcpl_1415));
  RMS_NORM_LOOP_1_1_and_15_nl <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), RMS_NORM_LOOP_1_1_mux1h_135_nl,
      RMS_NORM_LOOP_1_1_nor_seb);
  RMS_NORM_LOOP_1_1_mux1h_136_nl <= MUX1HOT_s_1_6_2((for_for_strm_in_tmp_sva_31_26(5)),
      attention_abs_qr_35_0_lpi_1_dfm_35, (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(35)),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(35)), (APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16(19)),
      attention_abs_4_qr_35_0_lpi_1_dfm_35, STD_LOGIC_VECTOR'( and_dcpl_1393 & and_dcpl_1398
      & RMS_NORM_LOOP_1_1_or_3_ssc & RMS_NORM_LOOP_1_1_or_1_ssc & and_dcpl_1415 &
      and_dcpl_1431));
  RMS_NORM_LOOP_1_1_mux1h_137_nl <= MUX1HOT_v_6_6_2(STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(for_for_strm_in_tmp_sva_31_26(5),
      1),6)), (attention_abs_qr_35_0_lpi_1_dfm_34_0(34 DOWNTO 29)), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(34
      DOWNTO 29)), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(34
      DOWNTO 29)), (APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16(18 DOWNTO 13)),
      (attention_abs_4_qr_35_0_lpi_1_dfm_34_0(34 DOWNTO 29)), STD_LOGIC_VECTOR'(
      and_dcpl_1393 & and_dcpl_1398 & RMS_NORM_LOOP_1_1_or_3_ssc & RMS_NORM_LOOP_1_1_or_1_ssc
      & and_dcpl_1415 & and_dcpl_1431));
  RMS_NORM_LOOP_1_1_mux1h_138_nl <= MUX1HOT_v_5_6_2((for_for_strm_in_tmp_sva_31_26(4
      DOWNTO 0)), (attention_abs_qr_35_0_lpi_1_dfm_34_0(28 DOWNTO 24)), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(28
      DOWNTO 24)), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(28
      DOWNTO 24)), (APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16(12 DOWNTO 8)), (attention_abs_4_qr_35_0_lpi_1_dfm_34_0(28
      DOWNTO 24)), STD_LOGIC_VECTOR'( and_dcpl_1393 & and_dcpl_1398 & RMS_NORM_LOOP_1_1_or_3_ssc
      & RMS_NORM_LOOP_1_1_or_1_ssc & and_dcpl_1415 & and_dcpl_1431));
  RMS_NORM_LOOP_1_1_mux1h_139_nl <= MUX1HOT_v_8_6_2((for_for_strm_in_tmp_sva_25_2(23
      DOWNTO 16)), (attention_abs_qr_35_0_lpi_1_dfm_34_0(23 DOWNTO 16)), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(23
      DOWNTO 16)), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(23
      DOWNTO 16)), (APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16(7 DOWNTO 0)), (attention_abs_4_qr_35_0_lpi_1_dfm_34_0(23
      DOWNTO 16)), STD_LOGIC_VECTOR'( and_dcpl_1393 & and_dcpl_1398 & RMS_NORM_LOOP_1_1_or_3_ssc
      & RMS_NORM_LOOP_1_1_or_1_ssc & and_dcpl_1415 & and_dcpl_1431));
  RMS_NORM_LOOP_1_1_mux1h_140_nl <= MUX1HOT_v_8_6_2((for_for_strm_in_tmp_sva_25_2(15
      DOWNTO 8)), (attention_abs_qr_35_0_lpi_1_dfm_34_0(15 DOWNTO 8)), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(15
      DOWNTO 8)), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(15 DOWNTO
      8)), reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd, (attention_abs_4_qr_35_0_lpi_1_dfm_34_0(15
      DOWNTO 8)), STD_LOGIC_VECTOR'( and_dcpl_1393 & and_dcpl_1398 & RMS_NORM_LOOP_1_1_or_3_ssc
      & RMS_NORM_LOOP_1_1_or_1_ssc & and_dcpl_1415 & and_dcpl_1431));
  RMS_NORM_LOOP_1_1_mux1h_141_nl <= MUX1HOT_v_8_6_2((for_for_strm_in_tmp_sva_25_2(7
      DOWNTO 0)), (attention_abs_qr_35_0_lpi_1_dfm_34_0(7 DOWNTO 0)), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(7
      DOWNTO 0)), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(7 DOWNTO
      0)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2 & reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0), (attention_abs_4_qr_35_0_lpi_1_dfm_34_0(7
      DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_1393 & and_dcpl_1398 & RMS_NORM_LOOP_1_1_or_3_ssc
      & RMS_NORM_LOOP_1_1_or_1_ssc & and_dcpl_1415 & and_dcpl_1431));
  RMS_NORM_LOOP_1_1_mux1h_142_nl <= MUX1HOT_s_1_6_2((for_for_strm_in_tmp_sva_31_26(5)),
      (operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_17_16(1)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(39)), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd(2)),
      QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39, (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(39)),
      STD_LOGIC_VECTOR'( and_dcpl_1393 & RMS_NORM_LOOP_1_1_or_4_itm & RMS_NORM_LOOP_1_1_or_2_ssc
      & and_dcpl_1415 & and_dcpl_1420 & and_dcpl_1436));
  RMS_NORM_LOOP_1_1_and_16_nl <= RMS_NORM_LOOP_1_1_mux1h_142_nl AND (NOT and_dcpl_1410)
      AND (NOT and_dcpl_1403);
  RMS_NORM_LOOP_1_1_mux1h_143_nl <= MUX1HOT_v_15_6_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(for_for_strm_in_tmp_sva_31_26),15)),
      STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_17_16(1),
      1),15)), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(38 DOWNTO 24)), STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd(2),
      1),15)), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(38 DOWNTO
      24)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(38 DOWNTO 24)), STD_LOGIC_VECTOR'(
      and_dcpl_1393 & RMS_NORM_LOOP_1_1_or_4_itm & RMS_NORM_LOOP_1_1_or_2_ssc & and_dcpl_1415
      & and_dcpl_1420 & and_dcpl_1436));
  RMS_NORM_LOOP_1_1_and_17_nl <= RMS_NORM_LOOP_1_1_mux1h_143_nl AND STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(NOT
      and_dcpl_1410, 1),15)) AND STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(NOT and_dcpl_1403,
      1),15));
  RMS_NORM_LOOP_1_1_mux1h_144_nl <= MUX1HOT_v_7_7_2((for_for_strm_in_tmp_sva_25_2(23
      DOWNTO 17)), STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_17_16(1),
      1),7)), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(23 DOWNTO 17)), STD_LOGIC_VECTOR'(
      "0000100"), STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd(2),
      1),7)), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(23 DOWNTO
      17)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(23 DOWNTO 17)), STD_LOGIC_VECTOR'(
      and_dcpl_1393 & RMS_NORM_LOOP_1_1_or_4_itm & RMS_NORM_LOOP_1_1_or_2_ssc & and_dcpl_1410
      & and_dcpl_1415 & and_dcpl_1420 & and_dcpl_1436));
  not_5114_nl <= NOT and_dcpl_1403;
  RMS_NORM_LOOP_1_1_and_18_nl <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), RMS_NORM_LOOP_1_1_mux1h_144_nl,
      not_5114_nl);
  RMS_NORM_LOOP_1_1_mux1h_145_nl <= MUX1HOT_s_1_6_2((for_for_strm_in_tmp_sva_25_2(16)),
      (operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_17_16(0)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(16)), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd(2)),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(16)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(16)),
      STD_LOGIC_VECTOR'( and_dcpl_1393 & RMS_NORM_LOOP_1_1_or_4_itm & RMS_NORM_LOOP_1_1_or_2_ssc
      & and_dcpl_1415 & and_dcpl_1420 & and_dcpl_1436));
  RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_3_nl <= NOT((NOT(RMS_NORM_LOOP_1_1_mux1h_145_nl
      OR and_dcpl_1410)) OR and_dcpl_1403);
  RMS_NORM_LOOP_1_1_mux1h_146_nl <= MUX1HOT_s_1_6_2((for_for_strm_in_tmp_sva_25_2(15)),
      operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_15,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(15)), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd(2)),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(15)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(15)),
      STD_LOGIC_VECTOR'( and_dcpl_1393 & RMS_NORM_LOOP_1_1_or_4_itm & RMS_NORM_LOOP_1_1_or_2_ssc
      & and_dcpl_1415 & and_dcpl_1420 & and_dcpl_1436));
  RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_4_nl <= NOT((NOT(RMS_NORM_LOOP_1_1_mux1h_146_nl
      OR and_dcpl_1410)) OR and_dcpl_1403);
  RMS_NORM_LOOP_1_1_mux1h_147_nl <= MUX1HOT_v_2_6_2((for_for_strm_in_tmp_sva_25_2(14
      DOWNTO 13)), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd(2
      DOWNTO 1)), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(14 DOWNTO 13)), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd(1
      DOWNTO 0)), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(14 DOWNTO
      13)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(14 DOWNTO 13)), STD_LOGIC_VECTOR'(
      and_dcpl_1393 & RMS_NORM_LOOP_1_1_or_4_itm & RMS_NORM_LOOP_1_1_or_2_ssc & and_dcpl_1415
      & and_dcpl_1420 & and_dcpl_1436));
  RMS_NORM_LOOP_1_1_and_19_nl <= RMS_NORM_LOOP_1_1_mux1h_147_nl AND STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(NOT
      and_dcpl_1410, 1),2)) AND STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(NOT and_dcpl_1403,
      1),2));
  RMS_NORM_LOOP_1_1_mux1h_148_nl <= MUX1HOT_s_1_6_2((for_for_strm_in_tmp_sva_25_2(12)),
      (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd(0)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(12)), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1(2)),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(12)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(12)),
      STD_LOGIC_VECTOR'( and_dcpl_1393 & RMS_NORM_LOOP_1_1_or_4_itm & RMS_NORM_LOOP_1_1_or_2_ssc
      & and_dcpl_1415 & and_dcpl_1420 & and_dcpl_1436));
  RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_5_nl <= NOT((NOT(RMS_NORM_LOOP_1_1_mux1h_148_nl
      OR and_dcpl_1410)) OR and_dcpl_1403);
  RMS_NORM_LOOP_1_1_mux1h_149_nl <= MUX1HOT_v_2_7_2((for_for_strm_in_tmp_sva_25_2(11
      DOWNTO 10)), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1(2
      DOWNTO 1)), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(11 DOWNTO 10)), STD_LOGIC_VECTOR'(
      "01"), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1(1
      DOWNTO 0)), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(11 DOWNTO
      10)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(11 DOWNTO 10)), STD_LOGIC_VECTOR'(
      and_dcpl_1393 & RMS_NORM_LOOP_1_1_or_5_cse & RMS_NORM_LOOP_1_1_or_2_ssc & and_dcpl_1410
      & and_dcpl_1415 & and_dcpl_1420 & and_dcpl_1436));
  RMS_NORM_LOOP_1_1_mux1h_150_nl <= MUX1HOT_s_1_6_2((for_for_strm_in_tmp_sva_25_2(9)),
      (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1(0)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(9)), reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2,
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(9)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(9)),
      STD_LOGIC_VECTOR'( and_dcpl_1393 & RMS_NORM_LOOP_1_1_or_5_cse & RMS_NORM_LOOP_1_1_or_2_ssc
      & and_dcpl_1415 & and_dcpl_1420 & and_dcpl_1436));
  RMS_NORM_LOOP_1_1_and_20_nl <= RMS_NORM_LOOP_1_1_mux1h_150_nl AND (NOT and_dcpl_1410);
  RMS_NORM_LOOP_1_1_mux1h_151_nl <= MUX1HOT_s_1_6_2((for_for_strm_in_tmp_sva_25_2(8)),
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(8)), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3(7)),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(8)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(8)),
      STD_LOGIC_VECTOR'( and_dcpl_1393 & RMS_NORM_LOOP_1_1_or_5_cse & RMS_NORM_LOOP_1_1_or_2_ssc
      & and_dcpl_1415 & and_dcpl_1420 & and_dcpl_1436));
  RMS_NORM_LOOP_1_1_or_13_nl <= RMS_NORM_LOOP_1_1_mux1h_151_nl OR and_dcpl_1410;
  RMS_NORM_LOOP_1_1_mux1h_152_nl <= MUX1HOT_v_2_7_2((for_for_strm_in_tmp_sva_25_2(7
      DOWNTO 6)), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3(7
      DOWNTO 6)), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(7 DOWNTO 6)), STD_LOGIC_VECTOR'(
      "01"), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3(6
      DOWNTO 5)), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(7 DOWNTO
      6)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(7 DOWNTO 6)), STD_LOGIC_VECTOR'(
      and_dcpl_1393 & RMS_NORM_LOOP_1_1_or_5_cse & RMS_NORM_LOOP_1_1_or_2_ssc & and_dcpl_1410
      & and_dcpl_1415 & and_dcpl_1420 & and_dcpl_1436));
  RMS_NORM_LOOP_1_1_mux1h_153_nl <= MUX1HOT_s_1_5_2((for_for_strm_in_tmp_sva_25_2(5)),
      (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3(5)),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(5)), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(5)),
      (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(5)), STD_LOGIC_VECTOR'( and_dcpl_1393
      & RMS_NORM_LOOP_1_1_or_5_cse & RMS_NORM_LOOP_1_1_or_2_ssc & and_dcpl_1420 &
      and_dcpl_1436));
  RMS_NORM_LOOP_1_1_or_14_nl <= RMS_NORM_LOOP_1_1_mux1h_153_nl OR and_dcpl_1415 OR
      and_dcpl_1410;
  RMS_NORM_LOOP_1_1_or_15_nl <= and_dcpl_1398 OR and_dcpl_1403 OR and_dcpl_1415 OR
      and_dcpl_1431;
  RMS_NORM_LOOP_1_1_mux1h_154_nl <= MUX1HOT_v_5_6_2((for_for_strm_in_tmp_sva_25_2(4
      DOWNTO 0)), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3(4
      DOWNTO 0)), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm(4 DOWNTO 0)), STD_LOGIC_VECTOR'(
      "10001"), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0(4 DOWNTO
      0)), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva(4 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_1393 & RMS_NORM_LOOP_1_1_or_15_nl & RMS_NORM_LOOP_1_1_or_2_ssc & and_dcpl_1410
      & and_dcpl_1420 & and_dcpl_1436));
  z_out_10 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(RMS_NORM_LOOP_1_1_and_14_nl
      & RMS_NORM_LOOP_1_1_and_15_nl & RMS_NORM_LOOP_1_1_mux1h_136_nl & RMS_NORM_LOOP_1_1_mux1h_137_nl
      & RMS_NORM_LOOP_1_1_mux1h_138_nl & RMS_NORM_LOOP_1_1_mux1h_139_nl & RMS_NORM_LOOP_1_1_mux1h_140_nl
      & RMS_NORM_LOOP_1_1_mux1h_141_nl) * SIGNED(RMS_NORM_LOOP_1_1_and_16_nl & RMS_NORM_LOOP_1_1_and_17_nl
      & RMS_NORM_LOOP_1_1_and_18_nl & RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_3_nl
      & RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_4_nl & RMS_NORM_LOOP_1_1_and_19_nl
      & RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_5_nl & RMS_NORM_LOOP_1_1_mux1h_149_nl
      & RMS_NORM_LOOP_1_1_and_20_nl & RMS_NORM_LOOP_1_1_or_13_nl & RMS_NORM_LOOP_1_1_mux1h_152_nl
      & RMS_NORM_LOOP_1_1_or_14_nl & RMS_NORM_LOOP_1_1_mux1h_154_nl)), 64));
  TRANSPOSE_LAST_TWO_DIMS_LOOP_3_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_mux_2_nl <= MUX_s_1_2_2(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd,
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd, and_dcpl_1447);
  TRANSPOSE_LAST_TWO_DIMS_LOOP_3_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_mux_3_nl <= MUX_s_1_2_2(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1,
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1, and_dcpl_1447);
  z_out_11 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'(
      TRANSPOSE_LAST_TWO_DIMS_LOOP_3_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_mux_2_nl & TRANSPOSE_LAST_TWO_DIMS_LOOP_3_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_mux_3_nl),
      2), 3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1), 2), 3), 3));
  nor_1397_nl <= NOT((fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1398_nl <= NOT((fsm_output(1)) OR or_dcpl_959);
  and_2128_nl <= (fsm_output(1)) AND (fsm_output(4)) AND (fsm_output(8));
  mux_2303_nl <= MUX_s_1_2_2(nor_1398_nl, and_2128_nl, fsm_output(2));
  mux_2302_nl <= MUX_s_1_2_2(nor_1397_nl, mux_2303_nl, fsm_output(3));
  mux_2301_nl <= MUX_s_1_2_2(mux_2302_nl, nor_1044_cse, fsm_output(6));
  mux_2300_nl <= MUX_s_1_2_2(mux_2301_nl, nor_1045_cse, fsm_output(7));
  RMS_NORM_LOOP_2_2_or_1_nl <= (and_dcpl_381 AND CONV_SL_1_1(fsm_output(1 DOWNTO
      0)=STD_LOGIC_VECTOR'("01")) AND and_dcpl_198) OR (mux_2300_nl AND (fsm_output(0))
      AND (NOT (fsm_output(5))));
  RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_mux_1_nl <= MUX_v_4_2_2(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0,
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2), RMS_NORM_LOOP_2_2_or_1_nl);
  z_out_12 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_mux_1_nl),
      5) + UNSIGNED'( "00001"), 5));
  and_2129_nl <= (NOT (fsm_output(8))) AND (fsm_output(4)) AND (fsm_output(1)) AND
      (fsm_output(2)) AND (fsm_output(0)) AND (NOT (fsm_output(3))) AND (fsm_output(5))
      AND nor_973_cse;
  RMS_NORM_LOOP_2_2_mux_28_nl <= MUX_v_53_2_2((APPLY_ROTARY_POS_EMB_LOOP_6_mul_3_itm(52
      DOWNTO 0)), STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm(51
      DOWNTO 0)),53)), and_2129_nl);
  mul_3_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39
      & QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0) * SIGNED(RMS_NORM_LOOP_2_2_mux_28_nl)),
      72));
  z_out_13_71_28 <= mul_3_nl(71 DOWNTO 28);
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_21_nl <= MUX_v_2_2_2((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(2
      DOWNTO 1)), STD_LOGIC_VECTOR'( reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1), and_dcpl_1248);
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_22_nl <= MUX_s_1_2_2((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd(0)),
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd, and_dcpl_1248);
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_23_nl <= MUX_s_1_2_2(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1,
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1, and_dcpl_1248);
  z_out <= MUX_v_16_16_2(attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_15_0, attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_15_0,
      (apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_15_8 & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_7
      & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_6 & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_5
      & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_4 & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_3
      & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_2 & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_1
      & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_0), attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_15_0,
      attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_15_0, attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_15_0,
      attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_15_0, attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_15_0,
      attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_15_0, attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_15_0,
      attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_15_0, attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_15_0,
      attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_15_0, attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_15_0,
      attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_15_0, attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_15_0,
      operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_21_nl & operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_22_nl
      & operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_23_nl);
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_22_nl <= MUX_s_1_2_2(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd, and_dcpl_1261);
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_23_nl <= MUX_s_1_2_2(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1, and_dcpl_1261);
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_24_nl <= MUX_s_1_2_2((reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(1)),
      reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0, and_dcpl_1261);
  operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_25_nl <= MUX_s_1_2_2((reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0)),
      reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1, and_dcpl_1261);
  z_out_1 <= MUX_v_16_16_2(attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_15_0,
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0, (apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_8
      & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_7 & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_6
      & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_5 & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_4
      & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_3 & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_2
      & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_1 & apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_0),
      attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_15_0,
      STD_LOGIC_VECTOR'( operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_22_nl &
      operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_23_nl & operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_24_nl
      & operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_25_nl));
  RMS_NORM_LOOP_2_2_mux_29_nl <= MUX_v_3_2_2(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd,
      STD_LOGIC_VECTOR'( reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(1))), and_dcpl_1273);
  RMS_NORM_LOOP_2_2_mux_30_nl <= MUX_s_1_2_2(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1,
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2(0)), and_dcpl_1273);
  z_out_2 <= MUX_v_40_16_2(attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1,
      attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3, attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3,
      attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3, attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3,
      RMS_NORM_LOOP_2_2_mux_29_nl & RMS_NORM_LOOP_2_2_mux_30_nl);
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    dut
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY dut IS
  PORT(
    clk : IN STD_LOGIC;
    en : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    strm_in_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    strm_in_rsc_vld : IN STD_LOGIC;
    strm_in_rsc_rdy : OUT STD_LOGIC;
    strm_out_rsc_dat : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    strm_out_rsc_vld : OUT STD_LOGIC;
    strm_out_rsc_rdy : IN STD_LOGIC
  );
END dut;

ARCHITECTURE v1 OF dut IS
  -- Interconnect Declarations
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_q_d : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d : STD_LOGIC_VECTOR (5 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d : STD_LOGIC_VECTOR (5 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL rms_norm_16_div_cmp_a : STD_LOGIC_VECTOR (71 DOWNTO 0);
  SIGNAL rms_norm_16_div_cmp_b : STD_LOGIC_VECTOR (60 DOWNTO 0);
  SIGNAL rms_norm_16_div_cmp_z : STD_LOGIC_VECTOR (71 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsc_clken : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsc_q : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsc_re : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsc_radr : STD_LOGIC_VECTOR (5 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsc_we : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsc_d : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsc_wadr : STD_LOGIC_VECTOR (5 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsc_clken : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsc_q : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsc_re : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsc_radr : STD_LOGIC_VECTOR (5 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsc_we : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsc_d : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsc_wadr : STD_LOGIC_VECTOR (5 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsc_clken : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsc_q : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsc_re : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsc_radr : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsc_we : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsc_d : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsc_wadr : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_iff : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_iff : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_iff : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_iff : STD_LOGIC;
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_iff : STD_LOGIC;

  SIGNAL rms_norm_16_div_cmp_a_1 : STD_LOGIC_VECTOR (71 DOWNTO 0);
  SIGNAL rms_norm_16_div_cmp_b_1 : STD_LOGIC_VECTOR (60 DOWNTO 0);
  SIGNAL rms_norm_16_div_cmp_z_1 : STD_LOGIC_VECTOR (71 DOWNTO 0);

  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsc_comp_d : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsc_comp_q : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsc_comp_radr : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsc_comp_wadr : STD_LOGIC_VECTOR (5
      DOWNTO 0);

  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsc_comp_d : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsc_comp_q : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsc_comp_radr : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsc_comp_wadr : STD_LOGIC_VECTOR (5
      DOWNTO 0);

  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsc_comp_d : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsc_comp_q : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsc_comp_radr : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsc_comp_wadr : STD_LOGIC_VECTOR
      (5 DOWNTO 0);

  COMPONENT dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_14_6_40_48_1_48_40_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
      re : OUT STD_LOGIC;
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      re_d : IN STD_LOGIC;
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_q : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_radr : STD_LOGIC_VECTOR (5 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_d : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr : STD_LOGIC_VECTOR (5 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_q_d_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);

  COMPONENT dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_15_6_40_48_1_48_40_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
      re : OUT STD_LOGIC;
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      re_d : IN STD_LOGIC;
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsci_q : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsci_radr : STD_LOGIC_VECTOR (5 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsci_d : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr : STD_LOGIC_VECTOR (5 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d_1 : STD_LOGIC_VECTOR (39 DOWNTO
      0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);

  COMPONENT dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_16_6_40_48_1_48_40_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
      re : OUT STD_LOGIC;
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      re_d : IN STD_LOGIC;
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsci_q : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsci_d : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsci_d_d : STD_LOGIC_VECTOR (39
      DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d_1 : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d_1 : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d_1 : STD_LOGIC_VECTOR
      (5 DOWNTO 0);

  COMPONENT dut_core
    PORT(
      clk : IN STD_LOGIC;
      en : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      strm_in_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      strm_in_rsc_vld : IN STD_LOGIC;
      strm_in_rsc_rdy : OUT STD_LOGIC;
      strm_out_rsc_dat : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      strm_out_rsc_vld : OUT STD_LOGIC;
      strm_out_rsc_rdy : IN STD_LOGIC;
      attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d : OUT STD_LOGIC;
      attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d : OUT STD_LOGIC_VECTOR (39 DOWNTO
          0);
      attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d : OUT STD_LOGIC_VECTOR (5 DOWNTO
          0);
      attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d : OUT STD_LOGIC_VECTOR (5 DOWNTO
          0);
      attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d : OUT STD_LOGIC_VECTOR (39 DOWNTO
          0);
      attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d : IN STD_LOGIC_VECTOR (39 DOWNTO
          0);
      attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d : OUT STD_LOGIC_VECTOR (5 DOWNTO
          0);
      attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d : OUT STD_LOGIC_VECTOR (5 DOWNTO
          0);
      attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d : IN STD_LOGIC_VECTOR (39
          DOWNTO 0);
      attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d : OUT STD_LOGIC_VECTOR
          (5 DOWNTO 0);
      attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d : OUT STD_LOGIC_VECTOR
          (5 DOWNTO 0);
      rms_norm_16_div_cmp_a : OUT STD_LOGIC_VECTOR (71 DOWNTO 0);
      rms_norm_16_div_cmp_b : OUT STD_LOGIC_VECTOR (60 DOWNTO 0);
      rms_norm_16_div_cmp_z : IN STD_LOGIC_VECTOR (71 DOWNTO 0);
      attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_pff : OUT STD_LOGIC;
      attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_pff : OUT STD_LOGIC;
      attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_pff : OUT STD_LOGIC;
      attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_pff : OUT STD_LOGIC;
      attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_pff : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL dut_core_inst_strm_in_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL dut_core_inst_strm_out_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL dut_core_inst_attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL dut_core_inst_attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL dut_core_inst_attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL dut_core_inst_attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL dut_core_inst_attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL dut_core_inst_attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL dut_core_inst_attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL dut_core_inst_attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d : STD_LOGIC_VECTOR
      (39 DOWNTO 0);
  SIGNAL dut_core_inst_attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL dut_core_inst_attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL dut_core_inst_rms_norm_16_div_cmp_a : STD_LOGIC_VECTOR (71 DOWNTO 0);
  SIGNAL dut_core_inst_rms_norm_16_div_cmp_b : STD_LOGIC_VECTOR (60 DOWNTO 0);
  SIGNAL dut_core_inst_rms_norm_16_div_cmp_z : STD_LOGIC_VECTOR (71 DOWNTO 0);

BEGIN
  rms_norm_16_div_cmp : work.mgc_comps.mgc_div
    GENERIC MAP(
      width_a => 72,
      width_b => 61,
      signd => 1
      )
    PORT MAP(
      a => rms_norm_16_div_cmp_a_1,
      b => rms_norm_16_div_cmp_b_1,
      z => rms_norm_16_div_cmp_z_1
    );
  rms_norm_16_div_cmp_a_1 <= rms_norm_16_div_cmp_a;
  rms_norm_16_div_cmp_b_1 <= rms_norm_16_div_cmp_b;
  rms_norm_16_div_cmp_z <= rms_norm_16_div_cmp_z_1;

  attention_2_1_16_16_4_4_k_cache_upd_rsc_comp : work.block_1r1w_rbw_pkg.BLOCK_1R1W_RBW
    GENERIC MAP(
      addr_width => 6,
      data_width => 40,
      depth => 48,
      latency => 1,
      suppress_sim_read_addr_range_errs => 1
      )
    PORT MAP(
      clk => clk,
      clken => attention_2_1_16_16_4_4_k_cache_upd_rsc_clken,
      d => attention_2_1_16_16_4_4_k_cache_upd_rsc_comp_d,
      q => attention_2_1_16_16_4_4_k_cache_upd_rsc_comp_q,
      radr => attention_2_1_16_16_4_4_k_cache_upd_rsc_comp_radr,
      re => attention_2_1_16_16_4_4_k_cache_upd_rsc_re,
      wadr => attention_2_1_16_16_4_4_k_cache_upd_rsc_comp_wadr,
      we => attention_2_1_16_16_4_4_k_cache_upd_rsc_we
    );
  attention_2_1_16_16_4_4_k_cache_upd_rsc_comp_d <= attention_2_1_16_16_4_4_k_cache_upd_rsc_d;
  attention_2_1_16_16_4_4_k_cache_upd_rsc_q <= attention_2_1_16_16_4_4_k_cache_upd_rsc_comp_q;
  attention_2_1_16_16_4_4_k_cache_upd_rsc_comp_radr <= attention_2_1_16_16_4_4_k_cache_upd_rsc_radr;
  attention_2_1_16_16_4_4_k_cache_upd_rsc_comp_wadr <= attention_2_1_16_16_4_4_k_cache_upd_rsc_wadr;

  attention_2_1_16_16_4_4_v_cache_upd_rsc_comp : work.block_1r1w_rbw_pkg.BLOCK_1R1W_RBW
    GENERIC MAP(
      addr_width => 6,
      data_width => 40,
      depth => 48,
      latency => 1,
      suppress_sim_read_addr_range_errs => 1
      )
    PORT MAP(
      clk => clk,
      clken => attention_2_1_16_16_4_4_v_cache_upd_rsc_clken,
      d => attention_2_1_16_16_4_4_v_cache_upd_rsc_comp_d,
      q => attention_2_1_16_16_4_4_v_cache_upd_rsc_comp_q,
      radr => attention_2_1_16_16_4_4_v_cache_upd_rsc_comp_radr,
      re => attention_2_1_16_16_4_4_v_cache_upd_rsc_re,
      wadr => attention_2_1_16_16_4_4_v_cache_upd_rsc_comp_wadr,
      we => attention_2_1_16_16_4_4_v_cache_upd_rsc_we
    );
  attention_2_1_16_16_4_4_v_cache_upd_rsc_comp_d <= attention_2_1_16_16_4_4_v_cache_upd_rsc_d;
  attention_2_1_16_16_4_4_v_cache_upd_rsc_q <= attention_2_1_16_16_4_4_v_cache_upd_rsc_comp_q;
  attention_2_1_16_16_4_4_v_cache_upd_rsc_comp_radr <= attention_2_1_16_16_4_4_v_cache_upd_rsc_radr;
  attention_2_1_16_16_4_4_v_cache_upd_rsc_comp_wadr <= attention_2_1_16_16_4_4_v_cache_upd_rsc_wadr;

  attention_2_1_16_16_4_4_k_proj_transposed_rsc_comp : work.block_1r1w_rbw_pkg.BLOCK_1R1W_RBW
    GENERIC MAP(
      addr_width => 6,
      data_width => 40,
      depth => 48,
      latency => 1,
      suppress_sim_read_addr_range_errs => 1
      )
    PORT MAP(
      clk => clk,
      clken => attention_2_1_16_16_4_4_k_proj_transposed_rsc_clken,
      d => attention_2_1_16_16_4_4_k_proj_transposed_rsc_comp_d,
      q => attention_2_1_16_16_4_4_k_proj_transposed_rsc_comp_q,
      radr => attention_2_1_16_16_4_4_k_proj_transposed_rsc_comp_radr,
      re => attention_2_1_16_16_4_4_k_proj_transposed_rsc_re,
      wadr => attention_2_1_16_16_4_4_k_proj_transposed_rsc_comp_wadr,
      we => attention_2_1_16_16_4_4_k_proj_transposed_rsc_we
    );
  attention_2_1_16_16_4_4_k_proj_transposed_rsc_comp_d <= attention_2_1_16_16_4_4_k_proj_transposed_rsc_d;
  attention_2_1_16_16_4_4_k_proj_transposed_rsc_q <= attention_2_1_16_16_4_4_k_proj_transposed_rsc_comp_q;
  attention_2_1_16_16_4_4_k_proj_transposed_rsc_comp_radr <= attention_2_1_16_16_4_4_k_proj_transposed_rsc_radr;
  attention_2_1_16_16_4_4_k_proj_transposed_rsc_comp_wadr <= attention_2_1_16_16_4_4_k_proj_transposed_rsc_wadr;

  attention_2_1_16_16_4_4_k_cache_upd_rsci : dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_14_6_40_48_1_48_40_1_gen
    PORT MAP(
      clken => attention_2_1_16_16_4_4_k_cache_upd_rsc_clken,
      q => attention_2_1_16_16_4_4_k_cache_upd_rsci_q,
      re => attention_2_1_16_16_4_4_k_cache_upd_rsc_re,
      radr => attention_2_1_16_16_4_4_k_cache_upd_rsci_radr,
      we => attention_2_1_16_16_4_4_k_cache_upd_rsc_we,
      d => attention_2_1_16_16_4_4_k_cache_upd_rsci_d,
      wadr => attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr,
      clken_d => attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d,
      d_d => attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d_1,
      q_d => attention_2_1_16_16_4_4_k_cache_upd_rsci_q_d_1,
      radr_d => attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d_1,
      re_d => attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_iff,
      wadr_d => attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d_1,
      we_d => attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_iff
    );
  attention_2_1_16_16_4_4_k_cache_upd_rsci_q <= attention_2_1_16_16_4_4_k_cache_upd_rsc_q;
  attention_2_1_16_16_4_4_k_cache_upd_rsc_radr <= attention_2_1_16_16_4_4_k_cache_upd_rsci_radr;
  attention_2_1_16_16_4_4_k_cache_upd_rsc_d <= attention_2_1_16_16_4_4_k_cache_upd_rsci_d;
  attention_2_1_16_16_4_4_k_cache_upd_rsc_wadr <= attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr;
  attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d_1 <= attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d;
  attention_2_1_16_16_4_4_k_cache_upd_rsci_q_d <= attention_2_1_16_16_4_4_k_cache_upd_rsci_q_d_1;
  attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d_1 <= attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d;
  attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d_1 <= attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d;

  attention_2_1_16_16_4_4_v_cache_upd_rsci : dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_15_6_40_48_1_48_40_1_gen
    PORT MAP(
      clken => attention_2_1_16_16_4_4_v_cache_upd_rsc_clken,
      q => attention_2_1_16_16_4_4_v_cache_upd_rsci_q,
      re => attention_2_1_16_16_4_4_v_cache_upd_rsc_re,
      radr => attention_2_1_16_16_4_4_v_cache_upd_rsci_radr,
      we => attention_2_1_16_16_4_4_v_cache_upd_rsc_we,
      d => attention_2_1_16_16_4_4_v_cache_upd_rsci_d,
      wadr => attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr,
      clken_d => attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d,
      d_d => attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d_1,
      q_d => attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d_1,
      radr_d => attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d_1,
      re_d => attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_iff,
      wadr_d => attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d_1,
      we_d => attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_iff
    );
  attention_2_1_16_16_4_4_v_cache_upd_rsci_q <= attention_2_1_16_16_4_4_v_cache_upd_rsc_q;
  attention_2_1_16_16_4_4_v_cache_upd_rsc_radr <= attention_2_1_16_16_4_4_v_cache_upd_rsci_radr;
  attention_2_1_16_16_4_4_v_cache_upd_rsc_d <= attention_2_1_16_16_4_4_v_cache_upd_rsci_d;
  attention_2_1_16_16_4_4_v_cache_upd_rsc_wadr <= attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr;
  attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d_1 <= attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d;
  attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d <= attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d_1;
  attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d_1 <= attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d;
  attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d_1 <= attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d;

  attention_2_1_16_16_4_4_k_proj_transposed_rsci : dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_16_6_40_48_1_48_40_1_gen
    PORT MAP(
      clken => attention_2_1_16_16_4_4_k_proj_transposed_rsc_clken,
      q => attention_2_1_16_16_4_4_k_proj_transposed_rsci_q,
      re => attention_2_1_16_16_4_4_k_proj_transposed_rsc_re,
      radr => attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr,
      we => attention_2_1_16_16_4_4_k_proj_transposed_rsc_we,
      d => attention_2_1_16_16_4_4_k_proj_transposed_rsci_d,
      wadr => attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr,
      clken_d => attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d,
      d_d => attention_2_1_16_16_4_4_k_proj_transposed_rsci_d_d,
      q_d => attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d_1,
      radr_d => attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d_1,
      re_d => attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_iff,
      wadr_d => attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d_1,
      we_d => attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_iff
    );
  attention_2_1_16_16_4_4_k_proj_transposed_rsci_q <= attention_2_1_16_16_4_4_k_proj_transposed_rsc_q;
  attention_2_1_16_16_4_4_k_proj_transposed_rsc_radr <= attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr;
  attention_2_1_16_16_4_4_k_proj_transposed_rsc_d <= attention_2_1_16_16_4_4_k_proj_transposed_rsci_d;
  attention_2_1_16_16_4_4_k_proj_transposed_rsc_wadr <= attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr;
  attention_2_1_16_16_4_4_k_proj_transposed_rsci_d_d <= attention_2_1_16_16_4_4_k_cache_upd_rsci_q_d;
  attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d <= attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d_1;
  attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d_1 <= attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d;
  attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d_1 <= attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d;

  dut_core_inst : dut_core
    PORT MAP(
      clk => clk,
      en => en,
      rst => rst,
      strm_in_rsc_dat => dut_core_inst_strm_in_rsc_dat,
      strm_in_rsc_vld => strm_in_rsc_vld,
      strm_in_rsc_rdy => strm_in_rsc_rdy,
      strm_out_rsc_dat => dut_core_inst_strm_out_rsc_dat,
      strm_out_rsc_vld => strm_out_rsc_vld,
      strm_out_rsc_rdy => strm_out_rsc_rdy,
      attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d => attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d,
      attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d => dut_core_inst_attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d,
      attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d => dut_core_inst_attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d,
      attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d => dut_core_inst_attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d,
      attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d => dut_core_inst_attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d,
      attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d => dut_core_inst_attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d,
      attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d => dut_core_inst_attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d,
      attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d => dut_core_inst_attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d,
      attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d => dut_core_inst_attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d,
      attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d => dut_core_inst_attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d,
      attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d => dut_core_inst_attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d,
      rms_norm_16_div_cmp_a => dut_core_inst_rms_norm_16_div_cmp_a,
      rms_norm_16_div_cmp_b => dut_core_inst_rms_norm_16_div_cmp_b,
      rms_norm_16_div_cmp_z => dut_core_inst_rms_norm_16_div_cmp_z,
      attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_pff => attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_iff,
      attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_pff => attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_iff,
      attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_pff => attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_iff,
      attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_pff => attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_iff,
      attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_pff => attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_iff
    );
  dut_core_inst_strm_in_rsc_dat <= strm_in_rsc_dat;
  strm_out_rsc_dat <= dut_core_inst_strm_out_rsc_dat;
  attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d <= dut_core_inst_attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d;
  attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d <= dut_core_inst_attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d;
  attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d <= dut_core_inst_attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d;
  attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d <= dut_core_inst_attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d;
  dut_core_inst_attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d <= attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d;
  attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d <= dut_core_inst_attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d;
  attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d <= dut_core_inst_attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d;
  dut_core_inst_attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d <= attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d;
  attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d <= dut_core_inst_attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d;
  attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d <= dut_core_inst_attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d;
  rms_norm_16_div_cmp_a <= dut_core_inst_rms_norm_16_div_cmp_a;
  rms_norm_16_div_cmp_b <= dut_core_inst_rms_norm_16_div_cmp_b;
  dut_core_inst_rms_norm_16_div_cmp_z <= rms_norm_16_div_cmp_z;

END v1;



