
//------> /opt/siemens/catapult/2024.1_2-1117371/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  localparam stallOff = 0; 
  wire                  stall_ctrl;
  assign stall_ctrl = stallOff;

  assign idat = dat;
  assign rdy = irdy && !stall_ctrl;
  assign ivld = vld && !stall_ctrl;

endmodule


//------> /opt/siemens/catapult/2024.1_2-1117371/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  localparam stallOff = 0; 
  wire stall_ctrl;
  assign stall_ctrl = stallOff;

  assign dat = idat;
  assign irdy = rdy && !stall_ctrl;
  assign vld = ivld && !stall_ctrl;

endmodule



//------> /opt/siemens/catapult/2024.1_2-1117371/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.v 
module mgc_div(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_a-1:0] z;  
   reg  [width_a-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  div_s(a,b,z);
	else
          div_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/siemens/catapult/2024.1_2-1117371/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)
// suppress_sim_read_addr_range_errs:  0 - report errors  1 - suppress errors

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 ,
  parameter suppress_sim_read_addr_range_errs = 1 
  
)( clk,clken,d,q,radr,re,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input  re;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" , syn_ramstyle = "block" *)
  reg [data_width-1:0] mem [depth-1:0];
  integer j;
  initial for (j = 0; j < depth; j = j + 1) mem[j] = 0;
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr READ_ENABLE re
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg re_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
          re_reg <= re;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./rtl_dutmgc_rom_33_32_20_1.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1_2/1117371 Production Release
//  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
// 
//  Generated by:   dr655@ecelinux-16.ece.cornell.edu
//  Generated date: Thu Nov 28 19:53:51 2024
// ----------------------------------------------------------------------

// 
module dutmgc_rom_33_32_20_1 (addr, data_out
);
  input [4:0]addr ;
  output [19:0]data_out ;


  // Constants for ROM dimensions
  parameter n_width    = 20;
  parameter n_size     = 32;
  parameter n_numports = 1;
  parameter n_addr_w   = 5;
  parameter n_inreg    = 0;
  parameter n_outreg   = 0;

  // Declare storage for memory elements
  reg [19:0] mem [31:0];

  // Declare output registers
  reg [19:0] data_out_t;

  // Initialize ROM contents
  initial begin: rom_init_blk
    mem[0] <= 20'b11110101111110101010;
    mem[1] <= 20'b11111101011111000111;
    mem[2] <= 20'b00000011110011011111;
    mem[3] <= 20'b11111100010011000010;
    mem[4] <= 20'b00110011110001011010;
    mem[5] <= 20'b11101110100010111101;
    mem[6] <= 20'b11101110111100000110;
    mem[7] <= 20'b00010111100010110000;
    mem[8] <= 20'b00001000000001000100;
    mem[9] <= 20'b00000011101100111101;
    mem[10] <= 20'b00000111010101100101;
    mem[11] <= 20'b00000100111101011001;
    mem[12] <= 20'b00000001100000111110;
    mem[13] <= 20'b11100001110001110100;
    mem[14] <= 20'b11111100011000010101;
    mem[15] <= 20'b11110111011000101010;
    mem[16] <= 20'b11011000011011010001;
    mem[17] <= 20'b10110011011011110001;
    mem[18] <= 20'b11111011110000001111;
    mem[19] <= 20'b11110101110011110011;
    mem[20] <= 20'b00010011000101001101;
    mem[21] <= 20'b11010000000001000001;
    mem[22] <= 20'b11111010010111000001;
    mem[23] <= 20'b11011110110011011101;
    mem[24] <= 20'b11111111100011101111;
    mem[25] <= 20'b00001010110111101011;
    mem[26] <= 20'b11111110010101011110;
    mem[27] <= 20'b00000000111010101100;
    mem[28] <= 20'b11011111111101000101;
    mem[29] <= 20'b00010011100111010101;
    mem[30] <= 20'b00111111100001111001;
    mem[31] <= 20'b11111000000011110000;
  end


  // Combinational ROM read block
  always@(*)
  begin
    data_out_t <= mem[addr];
  end

  // Output register assignment
  assign data_out = data_out_t;

endmodule



//------> ./rtl_dutmgc_rom_34_64_8_1.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1_2/1117371 Production Release
//  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
// 
//  Generated by:   dr655@ecelinux-16.ece.cornell.edu
//  Generated date: Thu Nov 28 19:53:51 2024
// ----------------------------------------------------------------------

// 
module dutmgc_rom_34_64_8_1 (addr, data_out
);
  input [5:0]addr ;
  output [7:0]data_out ;


  // Constants for ROM dimensions
  parameter n_width    = 8;
  parameter n_size     = 64;
  parameter n_numports = 1;
  parameter n_addr_w   = 6;
  parameter n_inreg    = 0;
  parameter n_outreg   = 0;

  // Declare storage for memory elements
  reg [7:0] mem [63:0];

  // Declare output registers
  reg [7:0] data_out_t;

  // Initialize ROM contents
  initial begin: rom_init_blk
    mem[0] <= 8'b10010010;
    mem[1] <= 8'b00100101;
    mem[2] <= 8'b10100110;
    mem[3] <= 8'b01100001;
    mem[4] <= 8'b10100101;
    mem[5] <= 8'b00100000;
    mem[6] <= 8'b01100001;
    mem[7] <= 8'b00000100;
    mem[8] <= 8'b01010001;
    mem[9] <= 8'b00010100;
    mem[10] <= 8'b10100101;
    mem[11] <= 8'b01010101;
    mem[12] <= 8'b10001000;
    mem[13] <= 8'b10010110;
    mem[14] <= 8'b10100000;
    mem[15] <= 8'b00011010;
    mem[16] <= 8'b01001001;
    mem[17] <= 8'b10100010;
    mem[18] <= 8'b01011001;
    mem[19] <= 8'b10101010;
    mem[20] <= 8'b10100010;
    mem[21] <= 8'b10100110;
    mem[22] <= 8'b00100100;
    mem[23] <= 8'b10100100;
    mem[24] <= 8'b00100110;
    mem[25] <= 8'b10100010;
    mem[26] <= 8'b01000000;
    mem[27] <= 8'b00010100;
    mem[28] <= 8'b00101001;
    mem[29] <= 8'b10011001;
    mem[30] <= 8'b00000010;
    mem[31] <= 8'b01100010;
    mem[32] <= 8'b10000110;
    mem[33] <= 8'b01011010;
    mem[34] <= 8'b10000100;
    mem[35] <= 8'b01010000;
    mem[36] <= 8'b01101010;
    mem[37] <= 8'b01011000;
    mem[38] <= 8'b01000000;
    mem[39] <= 8'b00100001;
    mem[40] <= 8'b01101001;
    mem[41] <= 8'b01010110;
    mem[42] <= 8'b10100110;
    mem[43] <= 8'b01000000;
    mem[44] <= 8'b01010001;
    mem[45] <= 8'b01101001;
    mem[46] <= 8'b01100100;
    mem[47] <= 8'b00011001;
    mem[48] <= 8'b00000001;
    mem[49] <= 8'b10010100;
    mem[50] <= 8'b01101000;
    mem[51] <= 8'b00001001;
    mem[52] <= 8'b00010001;
    mem[53] <= 8'b00010000;
    mem[54] <= 8'b00100100;
    mem[55] <= 8'b10000000;
    mem[56] <= 8'b00000000;
    mem[57] <= 8'b00011010;
    mem[58] <= 8'b01010110;
    mem[59] <= 8'b00010101;
    mem[60] <= 8'b00001000;
    mem[61] <= 8'b00001010;
    mem[62] <= 8'b00101000;
    mem[63] <= 8'b00101010;
  end


  // Combinational ROM read block
  always@(*)
  begin
    data_out_t <= mem[addr];
  end

  // Output register assignment
  assign data_out = data_out_t;

endmodule



//------> ./rtl_dutmgc_rom_35_64_8_1.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1_2/1117371 Production Release
//  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
// 
//  Generated by:   dr655@ecelinux-16.ece.cornell.edu
//  Generated date: Thu Nov 28 19:53:51 2024
// ----------------------------------------------------------------------

// 
module dutmgc_rom_35_64_8_1 (addr, data_out
);
  input [5:0]addr ;
  output [7:0]data_out ;


  // Constants for ROM dimensions
  parameter n_width    = 8;
  parameter n_size     = 64;
  parameter n_numports = 1;
  parameter n_addr_w   = 6;
  parameter n_inreg    = 0;
  parameter n_outreg   = 0;

  // Declare storage for memory elements
  reg [7:0] mem [63:0];

  // Declare output registers
  reg [7:0] data_out_t;

  // Initialize ROM contents
  initial begin: rom_init_blk
    mem[0] <= 8'b10010110;
    mem[1] <= 8'b01101001;
    mem[2] <= 8'b10101000;
    mem[3] <= 8'b10100101;
    mem[4] <= 8'b10000110;
    mem[5] <= 8'b10100100;
    mem[6] <= 8'b10011001;
    mem[7] <= 8'b01100110;
    mem[8] <= 8'b10100101;
    mem[9] <= 8'b01010010;
    mem[10] <= 8'b00000010;
    mem[11] <= 8'b01010101;
    mem[12] <= 8'b00000010;
    mem[13] <= 8'b01010110;
    mem[14] <= 8'b01000010;
    mem[15] <= 8'b10010110;
    mem[16] <= 8'b00010110;
    mem[17] <= 8'b01010110;
    mem[18] <= 8'b00000101;
    mem[19] <= 8'b00011010;
    mem[20] <= 8'b01101000;
    mem[21] <= 8'b01010100;
    mem[22] <= 8'b00011010;
    mem[23] <= 8'b01010101;
    mem[24] <= 8'b10011010;
    mem[25] <= 8'b01100101;
    mem[26] <= 8'b00000101;
    mem[27] <= 8'b01010010;
    mem[28] <= 8'b10010001;
    mem[29] <= 8'b00010000;
    mem[30] <= 8'b01000101;
    mem[31] <= 8'b00010101;
    mem[32] <= 8'b00011000;
    mem[33] <= 8'b01010110;
    mem[34] <= 8'b00001001;
    mem[35] <= 8'b01000001;
    mem[36] <= 8'b01010110;
    mem[37] <= 8'b01001010;
    mem[38] <= 8'b01101001;
    mem[39] <= 8'b10000110;
    mem[40] <= 8'b10101010;
    mem[41] <= 8'b10000100;
    mem[42] <= 8'b10100110;
    mem[43] <= 8'b00011000;
    mem[44] <= 8'b01011001;
    mem[45] <= 8'b00100001;
    mem[46] <= 8'b10000100;
    mem[47] <= 8'b10011010;
    mem[48] <= 8'b10010110;
    mem[49] <= 8'b10101010;
    mem[50] <= 8'b01001000;
    mem[51] <= 8'b00100001;
    mem[52] <= 8'b01010001;
    mem[53] <= 8'b00101000;
    mem[54] <= 8'b01101000;
    mem[55] <= 8'b01001001;
    mem[56] <= 8'b10000110;
    mem[57] <= 8'b01001001;
    mem[58] <= 8'b10010110;
    mem[59] <= 8'b10100101;
    mem[60] <= 8'b10011000;
    mem[61] <= 8'b10000110;
    mem[62] <= 8'b10100101;
    mem[63] <= 8'b01000100;
  end


  // Combinational ROM read block
  always@(*)
  begin
    data_out_t <= mem[addr];
  end

  // Output register assignment
  assign data_out = data_out_t;

endmodule



//------> ./rtl_dutmgc_rom_36_960_15_1.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1_2/1117371 Production Release
//  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
// 
//  Generated by:   dr655@ecelinux-16.ece.cornell.edu
//  Generated date: Thu Nov 28 19:53:51 2024
// ----------------------------------------------------------------------

// 
module dutmgc_rom_36_960_15_1 (addr, data_out
);
  input [9:0]addr ;
  output [14:0]data_out ;


  // Constants for ROM dimensions
  parameter n_width    = 15;
  parameter n_size     = 960;
  parameter n_numports = 1;
  parameter n_addr_w   = 10;
  parameter n_inreg    = 0;
  parameter n_outreg   = 0;

  // Declare storage for memory elements
  reg [14:0] mem [959:0];

  // Declare output registers
  reg [14:0] data_out_t;

  // Initialize ROM contents
  initial begin: rom_init_blk
    mem[0] <= 15'b000000000000000;
    mem[1] <= 15'b000000000000000;
    mem[2] <= 15'b000000000000000;
    mem[3] <= 15'b000000000000000;
    mem[4] <= 15'b000000000000000;
    mem[5] <= 15'b000000000000000;
    mem[6] <= 15'b000000000000000;
    mem[7] <= 15'b000000000000000;
    mem[8] <= 15'b000000000000000;
    mem[9] <= 15'b000000000000000;
    mem[10] <= 15'b000000000000000;
    mem[11] <= 15'b000000000000000;
    mem[12] <= 15'b000000000000000;
    mem[13] <= 15'b000000000000000;
    mem[14] <= 15'b000000000000000;
    mem[15] <= 15'b000000000000000;
    mem[16] <= 15'b000000000000000;
    mem[17] <= 15'b000000000000000;
    mem[18] <= 15'b000000000000000;
    mem[19] <= 15'b000000000000000;
    mem[20] <= 15'b000000000000000;
    mem[21] <= 15'b000000000000000;
    mem[22] <= 15'b000000000000000;
    mem[23] <= 15'b000000000000000;
    mem[24] <= 15'b000000000000000;
    mem[25] <= 15'b000000000000000;
    mem[26] <= 15'b000000000000000;
    mem[27] <= 15'b000000000000000;
    mem[28] <= 15'b000000000000000;
    mem[29] <= 15'b000000000000000;
    mem[30] <= 15'b000000000000000;
    mem[31] <= 15'b000000000000000;
    mem[32] <= 15'b000000000000000;
    mem[33] <= 15'b000000000000000;
    mem[34] <= 15'b000000000000000;
    mem[35] <= 15'b000000000000000;
    mem[36] <= 15'b000000000000000;
    mem[37] <= 15'b000000000000000;
    mem[38] <= 15'b000000000000000;
    mem[39] <= 15'b000000000000000;
    mem[40] <= 15'b000000000000000;
    mem[41] <= 15'b000000000000000;
    mem[42] <= 15'b000000000000000;
    mem[43] <= 15'b000000000000000;
    mem[44] <= 15'b000000000000000;
    mem[45] <= 15'b000000000000000;
    mem[46] <= 15'b000000000000000;
    mem[47] <= 15'b000000000000000;
    mem[48] <= 15'b000000000000000;
    mem[49] <= 15'b000000000000000;
    mem[50] <= 15'b000000000000000;
    mem[51] <= 15'b000000000000000;
    mem[52] <= 15'b000000000000000;
    mem[53] <= 15'b000000000000000;
    mem[54] <= 15'b000000000000000;
    mem[55] <= 15'b000000000000000;
    mem[56] <= 15'b000000000000000;
    mem[57] <= 15'b000000000000000;
    mem[58] <= 15'b000000000000000;
    mem[59] <= 15'b000000000000000;
    mem[60] <= 15'b000000000000000;
    mem[61] <= 15'b000000000000000;
    mem[62] <= 15'b000000000000000;
    mem[63] <= 15'b000000000000000;
    mem[64] <= 15'b000000000000000;
    mem[65] <= 15'b000000000000000;
    mem[66] <= 15'b000000000000000;
    mem[67] <= 15'b000000000000000;
    mem[68] <= 15'b000000000000000;
    mem[69] <= 15'b000000000000000;
    mem[70] <= 15'b000000000000000;
    mem[71] <= 15'b000000000000000;
    mem[72] <= 15'b000000000000000;
    mem[73] <= 15'b000000000000000;
    mem[74] <= 15'b000000000000000;
    mem[75] <= 15'b000000000000000;
    mem[76] <= 15'b000000000000000;
    mem[77] <= 15'b000000000000000;
    mem[78] <= 15'b000000000000000;
    mem[79] <= 15'b000000000000000;
    mem[80] <= 15'b000000000000000;
    mem[81] <= 15'b000000000000000;
    mem[82] <= 15'b000000000000000;
    mem[83] <= 15'b000000000000000;
    mem[84] <= 15'b000000000000000;
    mem[85] <= 15'b000000000000000;
    mem[86] <= 15'b000000000000000;
    mem[87] <= 15'b000000000000000;
    mem[88] <= 15'b000000000000000;
    mem[89] <= 15'b000000000000000;
    mem[90] <= 15'b000000000000000;
    mem[91] <= 15'b000000000000000;
    mem[92] <= 15'b000000000000000;
    mem[93] <= 15'b000000000000000;
    mem[94] <= 15'b000000000000000;
    mem[95] <= 15'b000000000000000;
    mem[96] <= 15'b100010100110001;
    mem[97] <= 15'b101011011001100;
    mem[98] <= 15'b110001101111111;
    mem[99] <= 15'b110110001001110;
    mem[100] <= 15'b111001001101011;
    mem[101] <= 15'b111011010110010;
    mem[102] <= 15'b111100110101111;
    mem[103] <= 15'b111101110110100;
    mem[104] <= 15'b111110100010100;
    mem[105] <= 15'b111110111110110;
    mem[106] <= 15'b111111010011111;
    mem[107] <= 15'b111111100011111;
    mem[108] <= 15'b111111101011000;
    mem[109] <= 15'b111111110000000;
    mem[110] <= 15'b111111110101000;
    mem[111] <= 15'b111111111011000;
    mem[112] <= 15'b111111111011001;
    mem[113] <= 15'b111111111101111;
    mem[114] <= 15'b111111111111111;
    mem[115] <= 15'b111111111101001;
    mem[116] <= 15'b111111111110000;
    mem[117] <= 15'b111111111110101;
    mem[118] <= 15'b111111111111000;
    mem[119] <= 15'b111111111111011;
    mem[120] <= 15'b111111111111100;
    mem[121] <= 15'b111111111111101;
    mem[122] <= 15'b111111111111110;
    mem[123] <= 15'b111111111111110;
    mem[124] <= 15'b111111111111111;
    mem[125] <= 15'b111111111111111;
    mem[126] <= 15'b111111111111111;
    mem[127] <= 15'b111111111111111;
    mem[128] <= 15'b111111111111111;
    mem[129] <= 15'b111111111111111;
    mem[130] <= 15'b111111111111111;
    mem[131] <= 15'b111111111111111;
    mem[132] <= 15'b111111111111111;
    mem[133] <= 15'b111111111111111;
    mem[134] <= 15'b111111111111111;
    mem[135] <= 15'b111111111111111;
    mem[136] <= 15'b111111111111111;
    mem[137] <= 15'b111111111111111;
    mem[138] <= 15'b111111111111111;
    mem[139] <= 15'b111111111111111;
    mem[140] <= 15'b000000000000000;
    mem[141] <= 15'b000000000000000;
    mem[142] <= 15'b000000000000000;
    mem[143] <= 15'b000000000000000;
    mem[144] <= 15'b100010100110001;
    mem[145] <= 15'b101011011001100;
    mem[146] <= 15'b110001101111111;
    mem[147] <= 15'b110110001001110;
    mem[148] <= 15'b111001001101011;
    mem[149] <= 15'b111011010110010;
    mem[150] <= 15'b111100110101111;
    mem[151] <= 15'b111101110110100;
    mem[152] <= 15'b111110100010100;
    mem[153] <= 15'b111110111110110;
    mem[154] <= 15'b111111010011111;
    mem[155] <= 15'b111111100011111;
    mem[156] <= 15'b111111101011000;
    mem[157] <= 15'b111111110000000;
    mem[158] <= 15'b111111110101000;
    mem[159] <= 15'b111111111011000;
    mem[160] <= 15'b111111111011001;
    mem[161] <= 15'b111111111101111;
    mem[162] <= 15'b111111111111111;
    mem[163] <= 15'b111111111101001;
    mem[164] <= 15'b111111111110000;
    mem[165] <= 15'b111111111110101;
    mem[166] <= 15'b111111111111000;
    mem[167] <= 15'b111111111111011;
    mem[168] <= 15'b111111111111100;
    mem[169] <= 15'b111111111111101;
    mem[170] <= 15'b111111111111110;
    mem[171] <= 15'b111111111111110;
    mem[172] <= 15'b111111111111111;
    mem[173] <= 15'b111111111111111;
    mem[174] <= 15'b111111111111111;
    mem[175] <= 15'b111111111111111;
    mem[176] <= 15'b111111111111111;
    mem[177] <= 15'b111111111111111;
    mem[178] <= 15'b111111111111111;
    mem[179] <= 15'b111111111111111;
    mem[180] <= 15'b111111111111111;
    mem[181] <= 15'b111111111111111;
    mem[182] <= 15'b111111111111111;
    mem[183] <= 15'b111111111111111;
    mem[184] <= 15'b111111111111111;
    mem[185] <= 15'b111111111111111;
    mem[186] <= 15'b111111111111111;
    mem[187] <= 15'b111111111111111;
    mem[188] <= 15'b000000000000000;
    mem[189] <= 15'b000000000000000;
    mem[190] <= 15'b000000000000000;
    mem[191] <= 15'b000000000000000;
    mem[192] <= 15'b100101010110111;
    mem[193] <= 15'b111010111000101;
    mem[194] <= 15'b001101001111100;
    mem[195] <= 15'b011011100100001;
    mem[196] <= 15'b100110010101000;
    mem[197] <= 15'b101110000111001;
    mem[198] <= 15'b110011101000001;
    mem[199] <= 15'b110111011101001;
    mem[200] <= 15'b111010001011001;
    mem[201] <= 15'b111011111111001;
    mem[202] <= 15'b111101010001110;
    mem[203] <= 15'b111110001000101;
    mem[204] <= 15'b111110101100110;
    mem[205] <= 15'b111111001000101;
    mem[206] <= 15'b111111011000000;
    mem[207] <= 15'b111111100100001;
    mem[208] <= 15'b111111101100101;
    mem[209] <= 15'b111111110011111;
    mem[210] <= 15'b111111110111101;
    mem[211] <= 15'b111111111000110;
    mem[212] <= 15'b111111111100011;
    mem[213] <= 15'b111111111110110;
    mem[214] <= 15'b111111111100011;
    mem[215] <= 15'b111111111101100;
    mem[216] <= 15'b111111111110010;
    mem[217] <= 15'b111111111110111;
    mem[218] <= 15'b111111111111001;
    mem[219] <= 15'b111111111111011;
    mem[220] <= 15'b111111111111101;
    mem[221] <= 15'b111111111111110;
    mem[222] <= 15'b111111111111110;
    mem[223] <= 15'b111111111111111;
    mem[224] <= 15'b111111111111111;
    mem[225] <= 15'b111111111111111;
    mem[226] <= 15'b111111111111111;
    mem[227] <= 15'b111111111111111;
    mem[228] <= 15'b111111111111111;
    mem[229] <= 15'b111111111111111;
    mem[230] <= 15'b111111111111111;
    mem[231] <= 15'b111111111111111;
    mem[232] <= 15'b111111111111111;
    mem[233] <= 15'b111111111111111;
    mem[234] <= 15'b111111111111111;
    mem[235] <= 15'b111111111111111;
    mem[236] <= 15'b111111111111111;
    mem[237] <= 15'b111111111111111;
    mem[238] <= 15'b111111111111111;
    mem[239] <= 15'b000000000000000;
    mem[240] <= 15'b100101010110111;
    mem[241] <= 15'b111010111000101;
    mem[242] <= 15'b001101001111100;
    mem[243] <= 15'b011011100100001;
    mem[244] <= 15'b100110010101000;
    mem[245] <= 15'b101110000111001;
    mem[246] <= 15'b110011101000001;
    mem[247] <= 15'b110111011101001;
    mem[248] <= 15'b111010001011001;
    mem[249] <= 15'b111011111111001;
    mem[250] <= 15'b111101010001110;
    mem[251] <= 15'b111110001000101;
    mem[252] <= 15'b111110101100110;
    mem[253] <= 15'b111111001000101;
    mem[254] <= 15'b111111011000000;
    mem[255] <= 15'b111111100100001;
    mem[256] <= 15'b111111101100101;
    mem[257] <= 15'b111111110011111;
    mem[258] <= 15'b111111110111101;
    mem[259] <= 15'b111111111000110;
    mem[260] <= 15'b111111111100011;
    mem[261] <= 15'b111111111110110;
    mem[262] <= 15'b111111111100011;
    mem[263] <= 15'b111111111101100;
    mem[264] <= 15'b111111111110010;
    mem[265] <= 15'b111111111110111;
    mem[266] <= 15'b111111111111001;
    mem[267] <= 15'b111111111111011;
    mem[268] <= 15'b111111111111101;
    mem[269] <= 15'b111111111111110;
    mem[270] <= 15'b111111111111110;
    mem[271] <= 15'b111111111111111;
    mem[272] <= 15'b111111111111111;
    mem[273] <= 15'b111111111111111;
    mem[274] <= 15'b111111111111111;
    mem[275] <= 15'b111111111111111;
    mem[276] <= 15'b111111111111111;
    mem[277] <= 15'b111111111111111;
    mem[278] <= 15'b111111111111111;
    mem[279] <= 15'b111111111111111;
    mem[280] <= 15'b111111111111111;
    mem[281] <= 15'b111111111111111;
    mem[282] <= 15'b111111111111111;
    mem[283] <= 15'b111111111111111;
    mem[284] <= 15'b111111111111111;
    mem[285] <= 15'b111111111111111;
    mem[286] <= 15'b111111111111111;
    mem[287] <= 15'b000000000000000;
    mem[288] <= 15'b000000101001111;
    mem[289] <= 15'b001101101010101;
    mem[290] <= 15'b100010110110100;
    mem[291] <= 15'b111000100010001;
    mem[292] <= 15'b001011010110001;
    mem[293] <= 15'b011010001100100;
    mem[294] <= 15'b100101010011001;
    mem[295] <= 15'b101101010110101;
    mem[296] <= 15'b110011000111100;
    mem[297] <= 15'b110111000101010;
    mem[298] <= 15'b111001111011000;
    mem[299] <= 15'b111011110100110;
    mem[300] <= 15'b111101001010010;
    mem[301] <= 15'b111110000010010;
    mem[302] <= 15'b111110101001100;
    mem[303] <= 15'b111111000111101;
    mem[304] <= 15'b111111011000101;
    mem[305] <= 15'b111111100101111;
    mem[306] <= 15'b111111101111001;
    mem[307] <= 15'b111111110010111;
    mem[308] <= 15'b111111110110111;
    mem[309] <= 15'b111111111000010;
    mem[310] <= 15'b111111111100000;
    mem[311] <= 15'b111111111110100;
    mem[312] <= 15'b111111111100010;
    mem[313] <= 15'b111111111101011;
    mem[314] <= 15'b111111111110010;
    mem[315] <= 15'b111111111110110;
    mem[316] <= 15'b111111111111001;
    mem[317] <= 15'b111111111111011;
    mem[318] <= 15'b111111111111101;
    mem[319] <= 15'b111111111111101;
    mem[320] <= 15'b111111111111110;
    mem[321] <= 15'b111111111111111;
    mem[322] <= 15'b111111111111111;
    mem[323] <= 15'b111111111111111;
    mem[324] <= 15'b111111111111111;
    mem[325] <= 15'b111111111111111;
    mem[326] <= 15'b111111111111111;
    mem[327] <= 15'b111111111111111;
    mem[328] <= 15'b111111111111111;
    mem[329] <= 15'b111111111111111;
    mem[330] <= 15'b111111111111111;
    mem[331] <= 15'b111111111111111;
    mem[332] <= 15'b111111111111111;
    mem[333] <= 15'b111111111111111;
    mem[334] <= 15'b111111111111111;
    mem[335] <= 15'b111111111111111;
    mem[336] <= 15'b000000101001111;
    mem[337] <= 15'b001101101010101;
    mem[338] <= 15'b100010110110100;
    mem[339] <= 15'b111000100010001;
    mem[340] <= 15'b001011010110001;
    mem[341] <= 15'b011010001100100;
    mem[342] <= 15'b100101010011001;
    mem[343] <= 15'b101101010110101;
    mem[344] <= 15'b110011000111100;
    mem[345] <= 15'b110111000101010;
    mem[346] <= 15'b111001111011000;
    mem[347] <= 15'b111011110100110;
    mem[348] <= 15'b111101001010010;
    mem[349] <= 15'b111110000010010;
    mem[350] <= 15'b111110101001100;
    mem[351] <= 15'b111111000111101;
    mem[352] <= 15'b111111011000101;
    mem[353] <= 15'b111111100101111;
    mem[354] <= 15'b111111101111001;
    mem[355] <= 15'b111111110010111;
    mem[356] <= 15'b111111110110111;
    mem[357] <= 15'b111111111000010;
    mem[358] <= 15'b111111111100000;
    mem[359] <= 15'b111111111110100;
    mem[360] <= 15'b111111111100010;
    mem[361] <= 15'b111111111101011;
    mem[362] <= 15'b111111111110010;
    mem[363] <= 15'b111111111110110;
    mem[364] <= 15'b111111111111001;
    mem[365] <= 15'b111111111111011;
    mem[366] <= 15'b111111111111101;
    mem[367] <= 15'b111111111111101;
    mem[368] <= 15'b111111111111110;
    mem[369] <= 15'b111111111111111;
    mem[370] <= 15'b111111111111111;
    mem[371] <= 15'b111111111111111;
    mem[372] <= 15'b111111111111111;
    mem[373] <= 15'b111111111111111;
    mem[374] <= 15'b111111111111111;
    mem[375] <= 15'b111111111111111;
    mem[376] <= 15'b111111111111111;
    mem[377] <= 15'b111111111111111;
    mem[378] <= 15'b111111111111111;
    mem[379] <= 15'b111111111111111;
    mem[380] <= 15'b111111111111111;
    mem[381] <= 15'b111111111111111;
    mem[382] <= 15'b111111111111111;
    mem[383] <= 15'b111111111111111;
    mem[384] <= 15'b010110001001010;
    mem[385] <= 15'b000000110011100;
    mem[386] <= 15'b000101011101111;
    mem[387] <= 15'b010111110010000;
    mem[388] <= 15'b101101111111101;
    mem[389] <= 15'b000010011111111;
    mem[390] <= 15'b010011010000111;
    mem[391] <= 15'b100000001011000;
    mem[392] <= 15'b101001101001011;
    mem[393] <= 15'b110000011100111;
    mem[394] <= 15'b110101010001000;
    mem[395] <= 15'b111000101000101;
    mem[396] <= 15'b111010111101101;
    mem[397] <= 15'b111100100001110;
    mem[398] <= 15'b111101101001110;
    mem[399] <= 15'b111110011001100;
    mem[400] <= 15'b111110111011001;
    mem[401] <= 15'b111111010000000;
    mem[402] <= 15'b111111011110100;
    mem[403] <= 15'b111111101011010;
    mem[404] <= 15'b111111110001100;
    mem[405] <= 15'b111111110111010;
    mem[406] <= 15'b111111111001111;
    mem[407] <= 15'b111111111010011;
    mem[408] <= 15'b111111111101011;
    mem[409] <= 15'b111111111111100;
    mem[410] <= 15'b111111111100111;
    mem[411] <= 15'b111111111101111;
    mem[412] <= 15'b111111111110100;
    mem[413] <= 15'b111111111111000;
    mem[414] <= 15'b111111111111010;
    mem[415] <= 15'b111111111111100;
    mem[416] <= 15'b111111111111101;
    mem[417] <= 15'b111111111111110;
    mem[418] <= 15'b111111111111110;
    mem[419] <= 15'b111111111111111;
    mem[420] <= 15'b111111111111111;
    mem[421] <= 15'b111111111111111;
    mem[422] <= 15'b111111111111111;
    mem[423] <= 15'b111111111111111;
    mem[424] <= 15'b111111111111111;
    mem[425] <= 15'b111111111111111;
    mem[426] <= 15'b111111111111111;
    mem[427] <= 15'b111111111111111;
    mem[428] <= 15'b111111111111111;
    mem[429] <= 15'b111111111111111;
    mem[430] <= 15'b111111111111111;
    mem[431] <= 15'b111111111111111;
    mem[432] <= 15'b010110001001010;
    mem[433] <= 15'b000000110011100;
    mem[434] <= 15'b000101011101111;
    mem[435] <= 15'b010111110010000;
    mem[436] <= 15'b101101111111101;
    mem[437] <= 15'b000010011111111;
    mem[438] <= 15'b010011010000111;
    mem[439] <= 15'b100000001011000;
    mem[440] <= 15'b101001101001011;
    mem[441] <= 15'b110000011100111;
    mem[442] <= 15'b110101010001000;
    mem[443] <= 15'b111000101000101;
    mem[444] <= 15'b111010111101101;
    mem[445] <= 15'b111100100001110;
    mem[446] <= 15'b111101101001110;
    mem[447] <= 15'b111110011001100;
    mem[448] <= 15'b111110111011001;
    mem[449] <= 15'b111111010000000;
    mem[450] <= 15'b111111011110100;
    mem[451] <= 15'b111111101011010;
    mem[452] <= 15'b111111110001100;
    mem[453] <= 15'b111111110111010;
    mem[454] <= 15'b111111111001111;
    mem[455] <= 15'b111111111010011;
    mem[456] <= 15'b111111111101011;
    mem[457] <= 15'b111111111111100;
    mem[458] <= 15'b111111111100111;
    mem[459] <= 15'b111111111101111;
    mem[460] <= 15'b111111111110100;
    mem[461] <= 15'b111111111111000;
    mem[462] <= 15'b111111111111010;
    mem[463] <= 15'b111111111111100;
    mem[464] <= 15'b111111111111101;
    mem[465] <= 15'b111111111111110;
    mem[466] <= 15'b111111111111110;
    mem[467] <= 15'b111111111111111;
    mem[468] <= 15'b111111111111111;
    mem[469] <= 15'b111111111111111;
    mem[470] <= 15'b111111111111111;
    mem[471] <= 15'b111111111111111;
    mem[472] <= 15'b111111111111111;
    mem[473] <= 15'b111111111111111;
    mem[474] <= 15'b111111111111111;
    mem[475] <= 15'b111111111111111;
    mem[476] <= 15'b111111111111111;
    mem[477] <= 15'b111111111111111;
    mem[478] <= 15'b111111111111111;
    mem[479] <= 15'b111111111111111;
    mem[480] <= 15'b010010001011110;
    mem[481] <= 15'b011100100110101;
    mem[482] <= 15'b000010001100001;
    mem[483] <= 15'b000011011011100;
    mem[484] <= 15'b010100011001011;
    mem[485] <= 15'b101010011001011;
    mem[486] <= 15'b111111010101111;
    mem[487] <= 15'b010000110100011;
    mem[488] <= 15'b011110010100110;
    mem[489] <= 15'b101000010100101;
    mem[490] <= 15'b101111100000100;
    mem[491] <= 15'b110100100110010;
    mem[492] <= 15'b111000001001101;
    mem[493] <= 15'b111010101000100;
    mem[494] <= 15'b111100010101011;
    mem[495] <= 15'b111101011110001;
    mem[496] <= 15'b111110010000010;
    mem[497] <= 15'b111110110110010;
    mem[498] <= 15'b111111001101110;
    mem[499] <= 15'b111111011110010;
    mem[500] <= 15'b111111101000100;
    mem[501] <= 15'b111111101111101;
    mem[502] <= 15'b111111110101111;
    mem[503] <= 15'b111111111000111;
    mem[504] <= 15'b111111111001110;
    mem[505] <= 15'b111111111101000;
    mem[506] <= 15'b111111111111001;
    mem[507] <= 15'b111111111100110;
    mem[508] <= 15'b111111111101110;
    mem[509] <= 15'b111111111110011;
    mem[510] <= 15'b111111111110111;
    mem[511] <= 15'b111111111111010;
    mem[512] <= 15'b111111111111100;
    mem[513] <= 15'b111111111111101;
    mem[514] <= 15'b111111111111110;
    mem[515] <= 15'b111111111111110;
    mem[516] <= 15'b111111111111111;
    mem[517] <= 15'b111111111111111;
    mem[518] <= 15'b111111111111111;
    mem[519] <= 15'b111111111111111;
    mem[520] <= 15'b111111111111111;
    mem[521] <= 15'b111111111111111;
    mem[522] <= 15'b111111111111111;
    mem[523] <= 15'b111111111111111;
    mem[524] <= 15'b111111111111111;
    mem[525] <= 15'b111111111111111;
    mem[526] <= 15'b111111111111111;
    mem[527] <= 15'b111111111111111;
    mem[528] <= 15'b010010001011110;
    mem[529] <= 15'b011100100110101;
    mem[530] <= 15'b000010001100001;
    mem[531] <= 15'b000011011011100;
    mem[532] <= 15'b010100011001011;
    mem[533] <= 15'b101010011001011;
    mem[534] <= 15'b111111010101111;
    mem[535] <= 15'b010000110100011;
    mem[536] <= 15'b011110010100110;
    mem[537] <= 15'b101000010100101;
    mem[538] <= 15'b101111100000100;
    mem[539] <= 15'b110100100110010;
    mem[540] <= 15'b111000001001101;
    mem[541] <= 15'b111010101000100;
    mem[542] <= 15'b111100010101011;
    mem[543] <= 15'b111101011110001;
    mem[544] <= 15'b111110010000010;
    mem[545] <= 15'b111110110110010;
    mem[546] <= 15'b111111001101110;
    mem[547] <= 15'b111111011110010;
    mem[548] <= 15'b111111101000100;
    mem[549] <= 15'b111111101111101;
    mem[550] <= 15'b111111110101111;
    mem[551] <= 15'b111111111000111;
    mem[552] <= 15'b111111111001110;
    mem[553] <= 15'b111111111101000;
    mem[554] <= 15'b111111111111001;
    mem[555] <= 15'b111111111100110;
    mem[556] <= 15'b111111111101110;
    mem[557] <= 15'b111111111110011;
    mem[558] <= 15'b111111111110111;
    mem[559] <= 15'b111111111111010;
    mem[560] <= 15'b111111111111100;
    mem[561] <= 15'b111111111111101;
    mem[562] <= 15'b111111111111110;
    mem[563] <= 15'b111111111111110;
    mem[564] <= 15'b111111111111111;
    mem[565] <= 15'b111111111111111;
    mem[566] <= 15'b111111111111111;
    mem[567] <= 15'b111111111111111;
    mem[568] <= 15'b111111111111111;
    mem[569] <= 15'b111111111111111;
    mem[570] <= 15'b111111111111111;
    mem[571] <= 15'b111111111111111;
    mem[572] <= 15'b111111111111111;
    mem[573] <= 15'b111111111111111;
    mem[574] <= 15'b111111111111111;
    mem[575] <= 15'b111111111111111;
    mem[576] <= 15'b111101011101101;
    mem[577] <= 15'b001111001001100;
    mem[578] <= 15'b011010100011101;
    mem[579] <= 15'b000001101110001;
    mem[580] <= 15'b000100000000010;
    mem[581] <= 15'b010101011100000;
    mem[582] <= 15'b101011011111000;
    mem[583] <= 15'b000000010011111;
    mem[584] <= 15'b010001100100101;
    mem[585] <= 15'b011110111001101;
    mem[586] <= 15'b101000110001001;
    mem[587] <= 15'b101111110101001;
    mem[588] <= 15'b110100110101110;
    mem[589] <= 15'b111000010100001;
    mem[590] <= 15'b111010101101010;
    mem[591] <= 15'b111100011001111;
    mem[592] <= 15'b111101100000010;
    mem[593] <= 15'b111110010100101;
    mem[594] <= 15'b111110110101000;
    mem[595] <= 15'b111111001111101;
    mem[596] <= 15'b111111011111101;
    mem[597] <= 15'b111111101001011;
    mem[598] <= 15'b111111110000001;
    mem[599] <= 15'b111111110110010;
    mem[600] <= 15'b111111111001010;
    mem[601] <= 15'b111111111001111;
    mem[602] <= 15'b111111111101001;
    mem[603] <= 15'b111111111111010;
    mem[604] <= 15'b111111111100110;
    mem[605] <= 15'b111111111101110;
    mem[606] <= 15'b111111111110100;
    mem[607] <= 15'b111111111110111;
    mem[608] <= 15'b111111111111010;
    mem[609] <= 15'b111111111111100;
    mem[610] <= 15'b111111111111101;
    mem[611] <= 15'b111111111111110;
    mem[612] <= 15'b111111111111110;
    mem[613] <= 15'b111111111111111;
    mem[614] <= 15'b111111111111111;
    mem[615] <= 15'b111111111111111;
    mem[616] <= 15'b111111111111111;
    mem[617] <= 15'b111111111111111;
    mem[618] <= 15'b111111111111111;
    mem[619] <= 15'b111111111111111;
    mem[620] <= 15'b111111111111111;
    mem[621] <= 15'b111111111111111;
    mem[622] <= 15'b111111111111111;
    mem[623] <= 15'b111111111111111;
    mem[624] <= 15'b111101011101101;
    mem[625] <= 15'b001111001001100;
    mem[626] <= 15'b011010100011101;
    mem[627] <= 15'b000001101110001;
    mem[628] <= 15'b000100000000010;
    mem[629] <= 15'b010101011100000;
    mem[630] <= 15'b101011011111000;
    mem[631] <= 15'b000000010011111;
    mem[632] <= 15'b010001100100101;
    mem[633] <= 15'b011110111001101;
    mem[634] <= 15'b101000110001001;
    mem[635] <= 15'b101111110101001;
    mem[636] <= 15'b110100110101110;
    mem[637] <= 15'b111000010100001;
    mem[638] <= 15'b111010101101010;
    mem[639] <= 15'b111100011001111;
    mem[640] <= 15'b111101100000010;
    mem[641] <= 15'b111110010100101;
    mem[642] <= 15'b111110110101000;
    mem[643] <= 15'b111111001111101;
    mem[644] <= 15'b111111011111101;
    mem[645] <= 15'b111111101001011;
    mem[646] <= 15'b111111110000001;
    mem[647] <= 15'b111111110110010;
    mem[648] <= 15'b111111111001010;
    mem[649] <= 15'b111111111001111;
    mem[650] <= 15'b111111111101001;
    mem[651] <= 15'b111111111111010;
    mem[652] <= 15'b111111111100110;
    mem[653] <= 15'b111111111101110;
    mem[654] <= 15'b111111111110100;
    mem[655] <= 15'b111111111110111;
    mem[656] <= 15'b111111111111010;
    mem[657] <= 15'b111111111111100;
    mem[658] <= 15'b111111111111101;
    mem[659] <= 15'b111111111111110;
    mem[660] <= 15'b111111111111110;
    mem[661] <= 15'b111111111111111;
    mem[662] <= 15'b111111111111111;
    mem[663] <= 15'b111111111111111;
    mem[664] <= 15'b111111111111111;
    mem[665] <= 15'b111111111111111;
    mem[666] <= 15'b111111111111111;
    mem[667] <= 15'b111111111111111;
    mem[668] <= 15'b111111111111111;
    mem[669] <= 15'b111111111111111;
    mem[670] <= 15'b111111111111111;
    mem[671] <= 15'b111111111111111;
    mem[672] <= 15'b110000001111111;
    mem[673] <= 15'b110111111110001;
    mem[674] <= 15'b000011100011110;
    mem[675] <= 15'b010011001100100;
    mem[676] <= 15'b000000010111000;
    mem[677] <= 15'b000110101000010;
    mem[678] <= 15'b011001101000011;
    mem[679] <= 15'b101111110000110;
    mem[680] <= 15'b000100000000101;
    mem[681] <= 15'b010100011101111;
    mem[682] <= 15'b100001000101101;
    mem[683] <= 15'b101010010110010;
    mem[684] <= 15'b110000111110011;
    mem[685] <= 15'b110101100110111;
    mem[686] <= 15'b111000110110010;
    mem[687] <= 15'b111011000101010;
    mem[688] <= 15'b111100101011010;
    mem[689] <= 15'b111101101111010;
    mem[690] <= 15'b111110011100001;
    mem[691] <= 15'b111110111011100;
    mem[692] <= 15'b111111010011000;
    mem[693] <= 15'b111111100000101;
    mem[694] <= 15'b111111101000110;
    mem[695] <= 15'b111111110010100;
    mem[696] <= 15'b111111110111111;
    mem[697] <= 15'b111111111010010;
    mem[698] <= 15'b111111111010101;
    mem[699] <= 15'b111111111101101;
    mem[700] <= 15'b111111111111101;
    mem[701] <= 15'b111111111101000;
    mem[702] <= 15'b111111111101111;
    mem[703] <= 15'b111111111110101;
    mem[704] <= 15'b111111111111000;
    mem[705] <= 15'b111111111111010;
    mem[706] <= 15'b111111111111100;
    mem[707] <= 15'b111111111111101;
    mem[708] <= 15'b111111111111110;
    mem[709] <= 15'b111111111111110;
    mem[710] <= 15'b111111111111111;
    mem[711] <= 15'b111111111111111;
    mem[712] <= 15'b111111111111111;
    mem[713] <= 15'b111111111111111;
    mem[714] <= 15'b111111111111111;
    mem[715] <= 15'b111111111111111;
    mem[716] <= 15'b111111111111111;
    mem[717] <= 15'b111111111111111;
    mem[718] <= 15'b111111111111111;
    mem[719] <= 15'b111111111111111;
    mem[720] <= 15'b110000001111111;
    mem[721] <= 15'b110111111110001;
    mem[722] <= 15'b000011100011110;
    mem[723] <= 15'b010011001100100;
    mem[724] <= 15'b000000010111000;
    mem[725] <= 15'b000110101000010;
    mem[726] <= 15'b011001101000011;
    mem[727] <= 15'b101111110000110;
    mem[728] <= 15'b000100000000101;
    mem[729] <= 15'b010100011101111;
    mem[730] <= 15'b100001000101101;
    mem[731] <= 15'b101010010110010;
    mem[732] <= 15'b110000111110011;
    mem[733] <= 15'b110101100110111;
    mem[734] <= 15'b111000110110010;
    mem[735] <= 15'b111011000101010;
    mem[736] <= 15'b111100101011010;
    mem[737] <= 15'b111101101111010;
    mem[738] <= 15'b111110011100001;
    mem[739] <= 15'b111110111011100;
    mem[740] <= 15'b111111010011000;
    mem[741] <= 15'b111111100000101;
    mem[742] <= 15'b111111101000110;
    mem[743] <= 15'b111111110010100;
    mem[744] <= 15'b111111110111111;
    mem[745] <= 15'b111111111010010;
    mem[746] <= 15'b111111111010101;
    mem[747] <= 15'b111111111101101;
    mem[748] <= 15'b111111111111101;
    mem[749] <= 15'b111111111101000;
    mem[750] <= 15'b111111111101111;
    mem[751] <= 15'b111111111110101;
    mem[752] <= 15'b111111111111000;
    mem[753] <= 15'b111111111111010;
    mem[754] <= 15'b111111111111100;
    mem[755] <= 15'b111111111111101;
    mem[756] <= 15'b111111111111110;
    mem[757] <= 15'b111111111111110;
    mem[758] <= 15'b111111111111111;
    mem[759] <= 15'b111111111111111;
    mem[760] <= 15'b111111111111111;
    mem[761] <= 15'b111111111111111;
    mem[762] <= 15'b111111111111111;
    mem[763] <= 15'b111111111111111;
    mem[764] <= 15'b111111111111111;
    mem[765] <= 15'b111111111111111;
    mem[766] <= 15'b111111111111111;
    mem[767] <= 15'b111111111111111;
    mem[768] <= 15'b110110101100000;
    mem[769] <= 15'b111100110000010;
    mem[770] <= 15'b101011000000100;
    mem[771] <= 15'b110010100001001;
    mem[772] <= 15'b001010001000111;
    mem[773] <= 15'b000000001100010;
    mem[774] <= 15'b001011101000001;
    mem[775] <= 15'b100000010110001;
    mem[776] <= 15'b110110010000110;
    mem[777] <= 15'b001001011011100;
    mem[778] <= 15'b011000101111001;
    mem[779] <= 15'b100100001100000;
    mem[780] <= 15'b101100100100100;
    mem[781] <= 15'b110010100010110;
    mem[782] <= 15'b110110101101100;
    mem[783] <= 15'b111001101000101;
    mem[784] <= 15'b111011101001101;
    mem[785] <= 15'b111101000010011;
    mem[786] <= 15'b111101111111010;
    mem[787] <= 15'b111110100101111;
    mem[788] <= 15'b111111000010100;
    mem[789] <= 15'b111111010101010;
    mem[790] <= 15'b111111100011100;
    mem[791] <= 15'b111111101101100;
    mem[792] <= 15'b111111110001110;
    mem[793] <= 15'b111111110110001;
    mem[794] <= 15'b111111111011110;
    mem[795] <= 15'b111111111011101;
    mem[796] <= 15'b111111111110010;
    mem[797] <= 15'b111111111100001;
    mem[798] <= 15'b111111111101011;
    mem[799] <= 15'b111111111110001;
    mem[800] <= 15'b111111111110110;
    mem[801] <= 15'b111111111111001;
    mem[802] <= 15'b111111111111011;
    mem[803] <= 15'b111111111111100;
    mem[804] <= 15'b111111111111101;
    mem[805] <= 15'b111111111111110;
    mem[806] <= 15'b111111111111111;
    mem[807] <= 15'b111111111111111;
    mem[808] <= 15'b111111111111111;
    mem[809] <= 15'b111111111111111;
    mem[810] <= 15'b111111111111111;
    mem[811] <= 15'b111111111111111;
    mem[812] <= 15'b111111111111111;
    mem[813] <= 15'b111111111111111;
    mem[814] <= 15'b111111111111111;
    mem[815] <= 15'b111111111111111;
    mem[816] <= 15'b110110101100000;
    mem[817] <= 15'b111100110000010;
    mem[818] <= 15'b101011000000100;
    mem[819] <= 15'b110010100001001;
    mem[820] <= 15'b001010001000111;
    mem[821] <= 15'b000000001100010;
    mem[822] <= 15'b001011101000001;
    mem[823] <= 15'b100000010110001;
    mem[824] <= 15'b110110010000110;
    mem[825] <= 15'b001001011011100;
    mem[826] <= 15'b011000101111001;
    mem[827] <= 15'b100100001100000;
    mem[828] <= 15'b101100100100100;
    mem[829] <= 15'b110010100010110;
    mem[830] <= 15'b110110101101100;
    mem[831] <= 15'b111001101000101;
    mem[832] <= 15'b111011101001101;
    mem[833] <= 15'b111101000010011;
    mem[834] <= 15'b111101111111010;
    mem[835] <= 15'b111110100101111;
    mem[836] <= 15'b111111000010100;
    mem[837] <= 15'b111111010101010;
    mem[838] <= 15'b111111100011100;
    mem[839] <= 15'b111111101101100;
    mem[840] <= 15'b111111110001110;
    mem[841] <= 15'b111111110110001;
    mem[842] <= 15'b111111111011110;
    mem[843] <= 15'b111111111011101;
    mem[844] <= 15'b111111111110010;
    mem[845] <= 15'b111111111100001;
    mem[846] <= 15'b111111111101011;
    mem[847] <= 15'b111111111110001;
    mem[848] <= 15'b111111111110110;
    mem[849] <= 15'b111111111111001;
    mem[850] <= 15'b111111111111011;
    mem[851] <= 15'b111111111111100;
    mem[852] <= 15'b111111111111101;
    mem[853] <= 15'b111111111111110;
    mem[854] <= 15'b111111111111111;
    mem[855] <= 15'b111111111111111;
    mem[856] <= 15'b111111111111111;
    mem[857] <= 15'b111111111111111;
    mem[858] <= 15'b111111111111111;
    mem[859] <= 15'b111111111111111;
    mem[860] <= 15'b111111111111111;
    mem[861] <= 15'b111111111111111;
    mem[862] <= 15'b111111111111111;
    mem[863] <= 15'b111111111111111;
    mem[864] <= 15'b000101101100000;
    mem[865] <= 15'b011010100010010;
    mem[866] <= 15'b111111010000100;
    mem[867] <= 15'b010101111101110;
    mem[868] <= 15'b011111010100101;
    mem[869] <= 15'b000010111100010;
    mem[870] <= 15'b000010110000100;
    mem[871] <= 15'b010011000101111;
    mem[872] <= 15'b101000111110101;
    mem[873] <= 15'b111110000111000;
    mem[874] <= 15'b001111110100101;
    mem[875] <= 15'b011101100101110;
    mem[876] <= 15'b100111110001101;
    mem[877] <= 15'b101111001010101;
    mem[878] <= 15'b110100010100010;
    mem[879] <= 15'b110111111100101;
    mem[880] <= 15'b111010011111100;
    mem[881] <= 15'b111100001110001;
    mem[882] <= 15'b111101011010100;
    mem[883] <= 15'b111110001110111;
    mem[884] <= 15'b111110110010011;
    mem[885] <= 15'b111111001011011;
    mem[886] <= 15'b111111011100100;
    mem[887] <= 15'b111111100111010;
    mem[888] <= 15'b111111101110110;
    mem[889] <= 15'b111111110101011;
    mem[890] <= 15'b111111111000100;
    mem[891] <= 15'b111111111001100;
    mem[892] <= 15'b111111111100110;
    mem[893] <= 15'b111111111111001;
    mem[894] <= 15'b111111111100101;
    mem[895] <= 15'b111111111101101;
    mem[896] <= 15'b111111111110011;
    mem[897] <= 15'b111111111110111;
    mem[898] <= 15'b111111111111010;
    mem[899] <= 15'b111111111111100;
    mem[900] <= 15'b111111111111101;
    mem[901] <= 15'b111111111111110;
    mem[902] <= 15'b111111111111110;
    mem[903] <= 15'b111111111111111;
    mem[904] <= 15'b111111111111111;
    mem[905] <= 15'b111111111111111;
    mem[906] <= 15'b111111111111111;
    mem[907] <= 15'b111111111111111;
    mem[908] <= 15'b111111111111111;
    mem[909] <= 15'b111111111111111;
    mem[910] <= 15'b111111111111111;
    mem[911] <= 15'b111111111111111;
    mem[912] <= 15'b000101101100000;
    mem[913] <= 15'b011010100010010;
    mem[914] <= 15'b111111010000100;
    mem[915] <= 15'b010101111101110;
    mem[916] <= 15'b011111010100101;
    mem[917] <= 15'b000010111100010;
    mem[918] <= 15'b000010110000100;
    mem[919] <= 15'b010011000101111;
    mem[920] <= 15'b101000111110101;
    mem[921] <= 15'b111110000111000;
    mem[922] <= 15'b001111110100101;
    mem[923] <= 15'b011101100101110;
    mem[924] <= 15'b100111110001101;
    mem[925] <= 15'b101111001010101;
    mem[926] <= 15'b110100010100010;
    mem[927] <= 15'b110111111100101;
    mem[928] <= 15'b111010011111100;
    mem[929] <= 15'b111100001110001;
    mem[930] <= 15'b111101011010100;
    mem[931] <= 15'b111110001110111;
    mem[932] <= 15'b111110110010011;
    mem[933] <= 15'b111111001011011;
    mem[934] <= 15'b111111011100100;
    mem[935] <= 15'b111111100111010;
    mem[936] <= 15'b111111101110110;
    mem[937] <= 15'b111111110101011;
    mem[938] <= 15'b111111111000100;
    mem[939] <= 15'b111111111001100;
    mem[940] <= 15'b111111111100110;
    mem[941] <= 15'b111111111111001;
    mem[942] <= 15'b111111111100101;
    mem[943] <= 15'b111111111101101;
    mem[944] <= 15'b111111111110011;
    mem[945] <= 15'b111111111110111;
    mem[946] <= 15'b111111111111010;
    mem[947] <= 15'b111111111111100;
    mem[948] <= 15'b111111111111101;
    mem[949] <= 15'b111111111111110;
    mem[950] <= 15'b111111111111110;
    mem[951] <= 15'b111111111111111;
    mem[952] <= 15'b111111111111111;
    mem[953] <= 15'b111111111111111;
    mem[954] <= 15'b111111111111111;
    mem[955] <= 15'b111111111111111;
    mem[956] <= 15'b111111111111111;
    mem[957] <= 15'b111111111111111;
    mem[958] <= 15'b111111111111111;
    mem[959] <= 15'b111111111111111;
  end


  // Combinational ROM read block
  always@(*)
  begin
    if ( addr >= 1'd0 && addr < 10'd960)
      data_out_t <= mem[addr];
    else
    begin
      data_out_t <= {(15){1'b0}};
    end
  end

  // Output register assignment
  assign data_out = data_out_t;

endmodule



//------> ./rtl_dutmgc_rom_37_960_13_1.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1_2/1117371 Production Release
//  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
// 
//  Generated by:   dr655@ecelinux-16.ece.cornell.edu
//  Generated date: Thu Nov 28 19:53:51 2024
// ----------------------------------------------------------------------

// 
module dutmgc_rom_37_960_13_1 (addr, data_out
);
  input [9:0]addr ;
  output [12:0]data_out ;


  // Constants for ROM dimensions
  parameter n_width    = 13;
  parameter n_size     = 960;
  parameter n_numports = 1;
  parameter n_addr_w   = 10;
  parameter n_inreg    = 0;
  parameter n_outreg   = 0;

  // Declare storage for memory elements
  reg [12:0] mem [959:0];

  // Declare output registers
  reg [12:0] data_out_t;

  // Initialize ROM contents
  initial begin: rom_init_blk
    mem[0] <= 13'b0000000000000;
    mem[1] <= 13'b0000000000000;
    mem[2] <= 13'b0000000000000;
    mem[3] <= 13'b0000000000000;
    mem[4] <= 13'b0000000000000;
    mem[5] <= 13'b0000000000000;
    mem[6] <= 13'b0000000000000;
    mem[7] <= 13'b0000000000000;
    mem[8] <= 13'b0000000000000;
    mem[9] <= 13'b0000000000000;
    mem[10] <= 13'b0000000000000;
    mem[11] <= 13'b0000000000000;
    mem[12] <= 13'b0000000000000;
    mem[13] <= 13'b0000000000000;
    mem[14] <= 13'b0000000000000;
    mem[15] <= 13'b0000000000000;
    mem[16] <= 13'b0000000000000;
    mem[17] <= 13'b0000000000000;
    mem[18] <= 13'b0000000000000;
    mem[19] <= 13'b0000000000000;
    mem[20] <= 13'b0000000000000;
    mem[21] <= 13'b0000000000000;
    mem[22] <= 13'b0000000000000;
    mem[23] <= 13'b0000000000000;
    mem[24] <= 13'b0000000000000;
    mem[25] <= 13'b0000000000000;
    mem[26] <= 13'b0000000000000;
    mem[27] <= 13'b0000000000000;
    mem[28] <= 13'b0000000000000;
    mem[29] <= 13'b0000000000000;
    mem[30] <= 13'b0000000000000;
    mem[31] <= 13'b0000000000000;
    mem[32] <= 13'b0000000000000;
    mem[33] <= 13'b0000000000000;
    mem[34] <= 13'b0000000000000;
    mem[35] <= 13'b0000000000000;
    mem[36] <= 13'b0000000000000;
    mem[37] <= 13'b0000000000000;
    mem[38] <= 13'b0000000000000;
    mem[39] <= 13'b0000000000000;
    mem[40] <= 13'b0000000000000;
    mem[41] <= 13'b0000000000000;
    mem[42] <= 13'b0000000000000;
    mem[43] <= 13'b0000000000000;
    mem[44] <= 13'b0000000000000;
    mem[45] <= 13'b0000000000000;
    mem[46] <= 13'b0000000000000;
    mem[47] <= 13'b0000000000000;
    mem[48] <= 13'b0000000000000;
    mem[49] <= 13'b0000000000000;
    mem[50] <= 13'b0000000000000;
    mem[51] <= 13'b0000000000000;
    mem[52] <= 13'b0000000000000;
    mem[53] <= 13'b0000000000000;
    mem[54] <= 13'b0000000000000;
    mem[55] <= 13'b0000000000000;
    mem[56] <= 13'b0000000000000;
    mem[57] <= 13'b0000000000000;
    mem[58] <= 13'b0000000000000;
    mem[59] <= 13'b0000000000000;
    mem[60] <= 13'b0000000000000;
    mem[61] <= 13'b0000000000000;
    mem[62] <= 13'b0000000000000;
    mem[63] <= 13'b0000000000000;
    mem[64] <= 13'b0000000000000;
    mem[65] <= 13'b0000000000000;
    mem[66] <= 13'b0000000000000;
    mem[67] <= 13'b0000000000000;
    mem[68] <= 13'b0000000000000;
    mem[69] <= 13'b0000000000000;
    mem[70] <= 13'b0000000000000;
    mem[71] <= 13'b0000000000000;
    mem[72] <= 13'b0000000000000;
    mem[73] <= 13'b0000000000000;
    mem[74] <= 13'b0000000000000;
    mem[75] <= 13'b0000000000000;
    mem[76] <= 13'b0000000000000;
    mem[77] <= 13'b0000000000000;
    mem[78] <= 13'b0000000000000;
    mem[79] <= 13'b0000000000000;
    mem[80] <= 13'b0000000000000;
    mem[81] <= 13'b0000000000000;
    mem[82] <= 13'b0000000000000;
    mem[83] <= 13'b0000000000000;
    mem[84] <= 13'b0000000000000;
    mem[85] <= 13'b0000000000000;
    mem[86] <= 13'b0000000000000;
    mem[87] <= 13'b0000000000000;
    mem[88] <= 13'b0000000000000;
    mem[89] <= 13'b0000000000000;
    mem[90] <= 13'b0000000000000;
    mem[91] <= 13'b0000000000000;
    mem[92] <= 13'b0000000000000;
    mem[93] <= 13'b0000000000000;
    mem[94] <= 13'b0000000000000;
    mem[95] <= 13'b0000000000000;
    mem[96] <= 13'b1011101101010;
    mem[97] <= 13'b1110000010100;
    mem[98] <= 13'b0000100110011;
    mem[99] <= 13'b0100010000110;
    mem[100] <= 13'b1001010010111;
    mem[101] <= 13'b1111110101110;
    mem[102] <= 13'b0111110011000;
    mem[103] <= 13'b0001000001110;
    mem[104] <= 13'b1011010111011;
    mem[105] <= 13'b0110101001010;
    mem[106] <= 13'b0010101101101;
    mem[107] <= 13'b1111011110000;
    mem[108] <= 13'b1100110001101;
    mem[109] <= 13'b1010100011001;
    mem[110] <= 13'b1000101101100;
    mem[111] <= 13'b0111001100100;
    mem[112] <= 13'b0101111100000;
    mem[113] <= 13'b0100111001101;
    mem[114] <= 13'b0100000010111;
    mem[115] <= 13'b0011010101110;
    mem[116] <= 13'b0010110000011;
    mem[117] <= 13'b0010010001100;
    mem[118] <= 13'b0001111000001;
    mem[119] <= 13'b0001100011001;
    mem[120] <= 13'b0001010001111;
    mem[121] <= 13'b0001000011100;
    mem[122] <= 13'b0000110111110;
    mem[123] <= 13'b0000101110000;
    mem[124] <= 13'b0000100110000;
    mem[125] <= 13'b0000011111011;
    mem[126] <= 13'b0000011001111;
    mem[127] <= 13'b0000010101010;
    mem[128] <= 13'b0000010001101;
    mem[129] <= 13'b0000001110100;
    mem[130] <= 13'b0000001100000;
    mem[131] <= 13'b0000001001111;
    mem[132] <= 13'b0000001000001;
    mem[133] <= 13'b0000000110110;
    mem[134] <= 13'b0000000101100;
    mem[135] <= 13'b0000000100100;
    mem[136] <= 13'b0000000011110;
    mem[137] <= 13'b0000000011001;
    mem[138] <= 13'b0000000010100;
    mem[139] <= 13'b0000000010001;
    mem[140] <= 13'b0000000001110;
    mem[141] <= 13'b0000000001011;
    mem[142] <= 13'b0000000001001;
    mem[143] <= 13'b0000000000111;
    mem[144] <= 13'b1011101101010;
    mem[145] <= 13'b1110000010100;
    mem[146] <= 13'b0000100110011;
    mem[147] <= 13'b0100010000110;
    mem[148] <= 13'b1001010010111;
    mem[149] <= 13'b1111110101110;
    mem[150] <= 13'b0111110011000;
    mem[151] <= 13'b0001000001110;
    mem[152] <= 13'b1011010111011;
    mem[153] <= 13'b0110101001010;
    mem[154] <= 13'b0010101101101;
    mem[155] <= 13'b1111011110000;
    mem[156] <= 13'b1100110001101;
    mem[157] <= 13'b1010100011001;
    mem[158] <= 13'b1000101101100;
    mem[159] <= 13'b0111001100100;
    mem[160] <= 13'b0101111100000;
    mem[161] <= 13'b0100111001101;
    mem[162] <= 13'b0100000010111;
    mem[163] <= 13'b0011010101110;
    mem[164] <= 13'b0010110000011;
    mem[165] <= 13'b0010010001100;
    mem[166] <= 13'b0001111000001;
    mem[167] <= 13'b0001100011001;
    mem[168] <= 13'b0001010001111;
    mem[169] <= 13'b0001000011100;
    mem[170] <= 13'b0000110111110;
    mem[171] <= 13'b0000101110000;
    mem[172] <= 13'b0000100110000;
    mem[173] <= 13'b0000011111011;
    mem[174] <= 13'b0000011001111;
    mem[175] <= 13'b0000010101010;
    mem[176] <= 13'b0000010001101;
    mem[177] <= 13'b0000001110100;
    mem[178] <= 13'b0000001100000;
    mem[179] <= 13'b0000001001111;
    mem[180] <= 13'b0000001000001;
    mem[181] <= 13'b0000000110110;
    mem[182] <= 13'b0000000101100;
    mem[183] <= 13'b0000000100100;
    mem[184] <= 13'b0000000011110;
    mem[185] <= 13'b0000000011001;
    mem[186] <= 13'b0000000010100;
    mem[187] <= 13'b0000000010001;
    mem[188] <= 13'b0000000001110;
    mem[189] <= 13'b0000000001011;
    mem[190] <= 13'b0000000001001;
    mem[191] <= 13'b0000000000111;
    mem[192] <= 13'b0100011000111;
    mem[193] <= 13'b1111100110000;
    mem[194] <= 13'b1101001110100;
    mem[195] <= 13'b0011011111011;
    mem[196] <= 13'b0110011110001;
    mem[197] <= 13'b1000101111110;
    mem[198] <= 13'b1011101001101;
    mem[199] <= 13'b1111110100011;
    mem[200] <= 13'b0101011101110;
    mem[201] <= 13'b1100100100111;
    mem[202] <= 13'b0101000001101;
    mem[203] <= 13'b1110101101101;
    mem[204] <= 13'b1001011011000;
    mem[205] <= 13'b0101000001110;
    mem[206] <= 13'b0001011000100;
    mem[207] <= 13'b1110010111100;
    mem[208] <= 13'b1011110111011;
    mem[209] <= 13'b1001110010111;
    mem[210] <= 13'b1000000101101;
    mem[211] <= 13'b0110101011100;
    mem[212] <= 13'b0101100000111;
    mem[213] <= 13'b0100100011001;
    mem[214] <= 13'b0011110000011;
    mem[215] <= 13'b0011000110011;
    mem[216] <= 13'b0010100011110;
    mem[217] <= 13'b0010000111001;
    mem[218] <= 13'b0001101111100;
    mem[219] <= 13'b0001011100000;
    mem[220] <= 13'b0001001100000;
    mem[221] <= 13'b0000111110110;
    mem[222] <= 13'b0000110011110;
    mem[223] <= 13'b0000101010101;
    mem[224] <= 13'b0000100011010;
    mem[225] <= 13'b0000011101001;
    mem[226] <= 13'b0000011000000;
    mem[227] <= 13'b0000010011110;
    mem[228] <= 13'b0000010000011;
    mem[229] <= 13'b0000001101100;
    mem[230] <= 13'b0000001011001;
    mem[231] <= 13'b0000001001001;
    mem[232] <= 13'b0000000111100;
    mem[233] <= 13'b0000000110010;
    mem[234] <= 13'b0000000101001;
    mem[235] <= 13'b0000000100010;
    mem[236] <= 13'b0000000011100;
    mem[237] <= 13'b0000000010111;
    mem[238] <= 13'b0000000010011;
    mem[239] <= 13'b0000000001111;
    mem[240] <= 13'b0100011000111;
    mem[241] <= 13'b1111100110000;
    mem[242] <= 13'b1101001110100;
    mem[243] <= 13'b0011011111011;
    mem[244] <= 13'b0110011110001;
    mem[245] <= 13'b1000101111110;
    mem[246] <= 13'b1011101001101;
    mem[247] <= 13'b1111110100011;
    mem[248] <= 13'b0101011101110;
    mem[249] <= 13'b1100100100111;
    mem[250] <= 13'b0101000001101;
    mem[251] <= 13'b1110101101101;
    mem[252] <= 13'b1001011011000;
    mem[253] <= 13'b0101000001110;
    mem[254] <= 13'b0001011000100;
    mem[255] <= 13'b1110010111100;
    mem[256] <= 13'b1011110111011;
    mem[257] <= 13'b1001110010111;
    mem[258] <= 13'b1000000101101;
    mem[259] <= 13'b0110101011100;
    mem[260] <= 13'b0101100000111;
    mem[261] <= 13'b0100100011001;
    mem[262] <= 13'b0011110000011;
    mem[263] <= 13'b0011000110011;
    mem[264] <= 13'b0010100011110;
    mem[265] <= 13'b0010000111001;
    mem[266] <= 13'b0001101111100;
    mem[267] <= 13'b0001011100000;
    mem[268] <= 13'b0001001100000;
    mem[269] <= 13'b0000111110110;
    mem[270] <= 13'b0000110011110;
    mem[271] <= 13'b0000101010101;
    mem[272] <= 13'b0000100011010;
    mem[273] <= 13'b0000011101001;
    mem[274] <= 13'b0000011000000;
    mem[275] <= 13'b0000010011110;
    mem[276] <= 13'b0000010000011;
    mem[277] <= 13'b0000001101100;
    mem[278] <= 13'b0000001011001;
    mem[279] <= 13'b0000001001001;
    mem[280] <= 13'b0000000111100;
    mem[281] <= 13'b0000000110010;
    mem[282] <= 13'b0000000101001;
    mem[283] <= 13'b0000000100010;
    mem[284] <= 13'b0000000011100;
    mem[285] <= 13'b0000000010111;
    mem[286] <= 13'b0000000010011;
    mem[287] <= 13'b0000000001111;
    mem[288] <= 13'b0010000100000;
    mem[289] <= 13'b1111000101011;
    mem[290] <= 13'b0001111101110;
    mem[291] <= 13'b1111001000010;
    mem[292] <= 13'b1101111101111;
    mem[293] <= 13'b0100110010100;
    mem[294] <= 13'b1000000000010;
    mem[295] <= 13'b1010010010011;
    mem[296] <= 13'b1101000101111;
    mem[297] <= 13'b0001000110100;
    mem[298] <= 13'b0110100010101;
    mem[299] <= 13'b1101100000010;
    mem[300] <= 13'b0101110100010;
    mem[301] <= 13'b1111010111010;
    mem[302] <= 13'b1001111110010;
    mem[303] <= 13'b0101011111101;
    mem[304] <= 13'b0001110001000;
    mem[305] <= 13'b1110101011001;
    mem[306] <= 13'b1100000111110;
    mem[307] <= 13'b1010000000111;
    mem[308] <= 13'b1000010001001;
    mem[309] <= 13'b0110110100101;
    mem[310] <= 13'b0101101000101;
    mem[311] <= 13'b0100101001101;
    mem[312] <= 13'b0011110101110;
    mem[313] <= 13'b0011001010110;
    mem[314] <= 13'b0010100111011;
    mem[315] <= 13'b0010001010001;
    mem[316] <= 13'b0001110010000;
    mem[317] <= 13'b0001011110001;
    mem[318] <= 13'b0001001101101;
    mem[319] <= 13'b0001000000000;
    mem[320] <= 13'b0000110100111;
    mem[321] <= 13'b0000101011101;
    mem[322] <= 13'b0000100100000;
    mem[323] <= 13'b0000011101110;
    mem[324] <= 13'b0000011000100;
    mem[325] <= 13'b0000010100010;
    mem[326] <= 13'b0000010000101;
    mem[327] <= 13'b0000001101110;
    mem[328] <= 13'b0000001011011;
    mem[329] <= 13'b0000001001011;
    mem[330] <= 13'b0000000111110;
    mem[331] <= 13'b0000000110011;
    mem[332] <= 13'b0000000101010;
    mem[333] <= 13'b0000000100010;
    mem[334] <= 13'b0000000011100;
    mem[335] <= 13'b0000000010111;
    mem[336] <= 13'b0010000100000;
    mem[337] <= 13'b1111000101011;
    mem[338] <= 13'b0001111101110;
    mem[339] <= 13'b1111001000010;
    mem[340] <= 13'b1101111101111;
    mem[341] <= 13'b0100110010100;
    mem[342] <= 13'b1000000000010;
    mem[343] <= 13'b1010010010011;
    mem[344] <= 13'b1101000101111;
    mem[345] <= 13'b0001000110100;
    mem[346] <= 13'b0110100010101;
    mem[347] <= 13'b1101100000010;
    mem[348] <= 13'b0101110100010;
    mem[349] <= 13'b1111010111010;
    mem[350] <= 13'b1001111110010;
    mem[351] <= 13'b0101011111101;
    mem[352] <= 13'b0001110001000;
    mem[353] <= 13'b1110101011001;
    mem[354] <= 13'b1100000111110;
    mem[355] <= 13'b1010000000111;
    mem[356] <= 13'b1000010001001;
    mem[357] <= 13'b0110110100101;
    mem[358] <= 13'b0101101000101;
    mem[359] <= 13'b0100101001101;
    mem[360] <= 13'b0011110101110;
    mem[361] <= 13'b0011001010110;
    mem[362] <= 13'b0010100111011;
    mem[363] <= 13'b0010001010001;
    mem[364] <= 13'b0001110010000;
    mem[365] <= 13'b0001011110001;
    mem[366] <= 13'b0001001101101;
    mem[367] <= 13'b0001000000000;
    mem[368] <= 13'b0000110100111;
    mem[369] <= 13'b0000101011101;
    mem[370] <= 13'b0000100100000;
    mem[371] <= 13'b0000011101110;
    mem[372] <= 13'b0000011000100;
    mem[373] <= 13'b0000010100010;
    mem[374] <= 13'b0000010000101;
    mem[375] <= 13'b0000001101110;
    mem[376] <= 13'b0000001011011;
    mem[377] <= 13'b0000001001011;
    mem[378] <= 13'b0000000111110;
    mem[379] <= 13'b0000000110011;
    mem[380] <= 13'b0000000101010;
    mem[381] <= 13'b0000000100010;
    mem[382] <= 13'b0000000011100;
    mem[383] <= 13'b0000000010111;
    mem[384] <= 13'b1111001000010;
    mem[385] <= 13'b1011101101011;
    mem[386] <= 13'b0011110101110;
    mem[387] <= 13'b0011100101111;
    mem[388] <= 13'b1010110100000;
    mem[389] <= 13'b1111111001111;
    mem[390] <= 13'b1010000011000;
    mem[391] <= 13'b1110101001000;
    mem[392] <= 13'b0001001001111;
    mem[393] <= 13'b0011100100101;
    mem[394] <= 13'b0110111000101;
    mem[395] <= 13'b1011101000011;
    mem[396] <= 13'b0001110101011;
    mem[397] <= 13'b1001011111001;
    mem[398] <= 13'b0010011100011;
    mem[399] <= 13'b1100100011011;
    mem[400] <= 13'b0111101000010;
    mem[401] <= 13'b0011100010000;
    mem[402] <= 13'b0000001001001;
    mem[403] <= 13'b1101010101111;
    mem[404] <= 13'b1011000001001;
    mem[405] <= 13'b1001000110000;
    mem[406] <= 13'b0111100000101;
    mem[407] <= 13'b0110001100110;
    mem[408] <= 13'b0101000111101;
    mem[409] <= 13'b0100001110011;
    mem[410] <= 13'b0011011111001;
    mem[411] <= 13'b0010111000001;
    mem[412] <= 13'b0010011000000;
    mem[413] <= 13'b0001111101100;
    mem[414] <= 13'b0001100111100;
    mem[415] <= 13'b0001010101011;
    mem[416] <= 13'b0001000110100;
    mem[417] <= 13'b0000111010010;
    mem[418] <= 13'b0000110000000;
    mem[419] <= 13'b0000100111101;
    mem[420] <= 13'b0000100000110;
    mem[421] <= 13'b0000011011000;
    mem[422] <= 13'b0000010110010;
    mem[423] <= 13'b0000010010011;
    mem[424] <= 13'b0000001111001;
    mem[425] <= 13'b0000001100100;
    mem[426] <= 13'b0000001010010;
    mem[427] <= 13'b0000001000100;
    mem[428] <= 13'b0000000111000;
    mem[429] <= 13'b0000000101110;
    mem[430] <= 13'b0000000100110;
    mem[431] <= 13'b0000000011111;
    mem[432] <= 13'b1111001000010;
    mem[433] <= 13'b1011101101011;
    mem[434] <= 13'b0011110101110;
    mem[435] <= 13'b0011100101111;
    mem[436] <= 13'b1010110100000;
    mem[437] <= 13'b1111111001111;
    mem[438] <= 13'b1010000011000;
    mem[439] <= 13'b1110101001000;
    mem[440] <= 13'b0001001001111;
    mem[441] <= 13'b0011100100101;
    mem[442] <= 13'b0110111000101;
    mem[443] <= 13'b1011101000011;
    mem[444] <= 13'b0001110101011;
    mem[445] <= 13'b1001011111001;
    mem[446] <= 13'b0010011100011;
    mem[447] <= 13'b1100100011011;
    mem[448] <= 13'b0111101000010;
    mem[449] <= 13'b0011100010000;
    mem[450] <= 13'b0000001001001;
    mem[451] <= 13'b1101010101111;
    mem[452] <= 13'b1011000001001;
    mem[453] <= 13'b1001000110000;
    mem[454] <= 13'b0111100000101;
    mem[455] <= 13'b0110001100110;
    mem[456] <= 13'b0101000111101;
    mem[457] <= 13'b0100001110011;
    mem[458] <= 13'b0011011111001;
    mem[459] <= 13'b0010111000001;
    mem[460] <= 13'b0010011000000;
    mem[461] <= 13'b0001111101100;
    mem[462] <= 13'b0001100111100;
    mem[463] <= 13'b0001010101011;
    mem[464] <= 13'b0001000110100;
    mem[465] <= 13'b0000111010010;
    mem[466] <= 13'b0000110000000;
    mem[467] <= 13'b0000100111101;
    mem[468] <= 13'b0000100000110;
    mem[469] <= 13'b0000011011000;
    mem[470] <= 13'b0000010110010;
    mem[471] <= 13'b0000010010011;
    mem[472] <= 13'b0000001111001;
    mem[473] <= 13'b0000001100100;
    mem[474] <= 13'b0000001010010;
    mem[475] <= 13'b0000001000100;
    mem[476] <= 13'b0000000111000;
    mem[477] <= 13'b0000000101110;
    mem[478] <= 13'b0000000100110;
    mem[479] <= 13'b0000000011111;
    mem[480] <= 13'b0101010000011;
    mem[481] <= 13'b0101011000101;
    mem[482] <= 13'b1110100101000;
    mem[483] <= 13'b1001010111100;
    mem[484] <= 13'b1101101011010;
    mem[485] <= 13'b1000011110101;
    mem[486] <= 13'b1111111111100;
    mem[487] <= 13'b1011100000001;
    mem[488] <= 13'b0000101110011;
    mem[489] <= 13'b0011011010000;
    mem[490] <= 13'b0101101101001;
    mem[491] <= 13'b1000111000100;
    mem[492] <= 13'b1101010110100;
    mem[493] <= 13'b0011010100111;
    mem[494] <= 13'b1010110000011;
    mem[495] <= 13'b0011100001100;
    mem[496] <= 13'b1101011100001;
    mem[497] <= 13'b1000010111001;
    mem[498] <= 13'b0100001001100;
    mem[499] <= 13'b0000101010010;
    mem[500] <= 13'b1101110000110;
    mem[501] <= 13'b1011010111001;
    mem[502] <= 13'b1001011000101;
    mem[503] <= 13'b0111101111111;
    mem[504] <= 13'b0110011001100;
    mem[505] <= 13'b0101010010000;
    mem[506] <= 13'b0100010111000;
    mem[507] <= 13'b0011100110010;
    mem[508] <= 13'b0010111110001;
    mem[509] <= 13'b0010011100111;
    mem[510] <= 13'b0010000001100;
    mem[511] <= 13'b0001101010110;
    mem[512] <= 13'b0001011000010;
    mem[513] <= 13'b0001001000110;
    mem[514] <= 13'b0000111100000;
    mem[515] <= 13'b0000110001100;
    mem[516] <= 13'b0000101000111;
    mem[517] <= 13'b0000100001110;
    mem[518] <= 13'b0000011011111;
    mem[519] <= 13'b0000010111000;
    mem[520] <= 13'b0000010011000;
    mem[521] <= 13'b0000001111101;
    mem[522] <= 13'b0000001100111;
    mem[523] <= 13'b0000001010101;
    mem[524] <= 13'b0000001000110;
    mem[525] <= 13'b0000000111010;
    mem[526] <= 13'b0000000110000;
    mem[527] <= 13'b0000000100111;
    mem[528] <= 13'b0101010000011;
    mem[529] <= 13'b0101011000101;
    mem[530] <= 13'b1110100101000;
    mem[531] <= 13'b1001010111100;
    mem[532] <= 13'b1101101011010;
    mem[533] <= 13'b1000011110101;
    mem[534] <= 13'b1111111111100;
    mem[535] <= 13'b1011100000001;
    mem[536] <= 13'b0000101110011;
    mem[537] <= 13'b0011011010000;
    mem[538] <= 13'b0101101101001;
    mem[539] <= 13'b1000111000100;
    mem[540] <= 13'b1101010110100;
    mem[541] <= 13'b0011010100111;
    mem[542] <= 13'b1010110000011;
    mem[543] <= 13'b0011100001100;
    mem[544] <= 13'b1101011100001;
    mem[545] <= 13'b1000010111001;
    mem[546] <= 13'b0100001001100;
    mem[547] <= 13'b0000101010010;
    mem[548] <= 13'b1101110000110;
    mem[549] <= 13'b1011010111001;
    mem[550] <= 13'b1001011000101;
    mem[551] <= 13'b0111101111111;
    mem[552] <= 13'b0110011001100;
    mem[553] <= 13'b0101010010000;
    mem[554] <= 13'b0100010111000;
    mem[555] <= 13'b0011100110010;
    mem[556] <= 13'b0010111110001;
    mem[557] <= 13'b0010011100111;
    mem[558] <= 13'b0010000001100;
    mem[559] <= 13'b0001101010110;
    mem[560] <= 13'b0001011000010;
    mem[561] <= 13'b0001001000110;
    mem[562] <= 13'b0000111100000;
    mem[563] <= 13'b0000110001100;
    mem[564] <= 13'b0000101000111;
    mem[565] <= 13'b0000100001110;
    mem[566] <= 13'b0000011011111;
    mem[567] <= 13'b0000010111000;
    mem[568] <= 13'b0000010011000;
    mem[569] <= 13'b0000001111101;
    mem[570] <= 13'b0000001100111;
    mem[571] <= 13'b0000001010101;
    mem[572] <= 13'b0000001000110;
    mem[573] <= 13'b0000000111010;
    mem[574] <= 13'b0000000110000;
    mem[575] <= 13'b0000000100111;
    mem[576] <= 13'b1100001111000;
    mem[577] <= 13'b0011101000011;
    mem[578] <= 13'b1000001110110;
    mem[579] <= 13'b0010011001001;
    mem[580] <= 13'b1100101110001;
    mem[581] <= 13'b1111100101110;
    mem[582] <= 13'b1001010000000;
    mem[583] <= 13'b1111111111111;
    mem[584] <= 13'b1011000101010;
    mem[585] <= 13'b0000000110101;
    mem[586] <= 13'b0010101011110;
    mem[587] <= 13'b0101000100001;
    mem[588] <= 13'b1000010000100;
    mem[589] <= 13'b1100110100010;
    mem[590] <= 13'b0010110111100;
    mem[591] <= 13'b1010011000010;
    mem[592] <= 13'b0011001100000;
    mem[593] <= 13'b1101001001111;
    mem[594] <= 13'b1000001000101;
    mem[595] <= 13'b0011111110000;
    mem[596] <= 13'b0000100000000;
    mem[597] <= 13'b1101101000000;
    mem[598] <= 13'b1011010000100;
    mem[599] <= 13'b1001010010111;
    mem[600] <= 13'b0111101011010;
    mem[601] <= 13'b0110010101100;
    mem[602] <= 13'b0101001110110;
    mem[603] <= 13'b0100010100010;
    mem[604] <= 13'b0011100100001;
    mem[605] <= 13'b0010111100010;
    mem[606] <= 13'b0010011011011;
    mem[607] <= 13'b0010000000001;
    mem[608] <= 13'b0001101001111;
    mem[609] <= 13'b0001010111011;
    mem[610] <= 13'b0001001000001;
    mem[611] <= 13'b0000111011100;
    mem[612] <= 13'b0000110001001;
    mem[613] <= 13'b0000101000100;
    mem[614] <= 13'b0000100001011;
    mem[615] <= 13'b0000011011101;
    mem[616] <= 13'b0000010110110;
    mem[617] <= 13'b0000010010110;
    mem[618] <= 13'b0000001111100;
    mem[619] <= 13'b0000001100110;
    mem[620] <= 13'b0000001010100;
    mem[621] <= 13'b0000001000101;
    mem[622] <= 13'b0000000111001;
    mem[623] <= 13'b0000000101111;
    mem[624] <= 13'b1100001111000;
    mem[625] <= 13'b0011101000011;
    mem[626] <= 13'b1000001110110;
    mem[627] <= 13'b0010011001001;
    mem[628] <= 13'b1100101110001;
    mem[629] <= 13'b1111100101110;
    mem[630] <= 13'b1001010000000;
    mem[631] <= 13'b1111111111111;
    mem[632] <= 13'b1011000101010;
    mem[633] <= 13'b0000000110101;
    mem[634] <= 13'b0010101011110;
    mem[635] <= 13'b0101000100001;
    mem[636] <= 13'b1000010000100;
    mem[637] <= 13'b1100110100010;
    mem[638] <= 13'b0010110111100;
    mem[639] <= 13'b1010011000010;
    mem[640] <= 13'b0011001100000;
    mem[641] <= 13'b1101001001111;
    mem[642] <= 13'b1000001000101;
    mem[643] <= 13'b0011111110000;
    mem[644] <= 13'b0000100000000;
    mem[645] <= 13'b1101101000000;
    mem[646] <= 13'b1011010000100;
    mem[647] <= 13'b1001010010111;
    mem[648] <= 13'b0111101011010;
    mem[649] <= 13'b0110010101100;
    mem[650] <= 13'b0101001110110;
    mem[651] <= 13'b0100010100010;
    mem[652] <= 13'b0011100100001;
    mem[653] <= 13'b0010111100010;
    mem[654] <= 13'b0010011011011;
    mem[655] <= 13'b0010000000001;
    mem[656] <= 13'b0001101001111;
    mem[657] <= 13'b0001010111011;
    mem[658] <= 13'b0001001000001;
    mem[659] <= 13'b0000111011100;
    mem[660] <= 13'b0000110001001;
    mem[661] <= 13'b0000101000100;
    mem[662] <= 13'b0000100001011;
    mem[663] <= 13'b0000011011101;
    mem[664] <= 13'b0000010110110;
    mem[665] <= 13'b0000010010110;
    mem[666] <= 13'b0000001111100;
    mem[667] <= 13'b0000001100110;
    mem[668] <= 13'b0000001010100;
    mem[669] <= 13'b0000001000101;
    mem[670] <= 13'b0000000111001;
    mem[671] <= 13'b0000000101111;
    mem[672] <= 13'b0100000110000;
    mem[673] <= 13'b0001110111100;
    mem[674] <= 13'b0000001100101;
    mem[675] <= 13'b0100100010110;
    mem[676] <= 13'b0010010011100;
    mem[677] <= 13'b1000110110010;
    mem[678] <= 13'b0110011111010;
    mem[679] <= 13'b1011110100110;
    mem[680] <= 13'b1111101111111;
    mem[681] <= 13'b1001010001000;
    mem[682] <= 13'b1101100010101;
    mem[683] <= 13'b0000000000000;
    mem[684] <= 13'b0010011100010;
    mem[685] <= 13'b0101111001001;
    mem[686] <= 13'b1010101111101;
    mem[687] <= 13'b0001000110100;
    mem[688] <= 13'b1000110111001;
    mem[689] <= 13'b0001111010000;
    mem[690] <= 13'b1100000110001;
    mem[691] <= 13'b0111010000110;
    mem[692] <= 13'b0011001110110;
    mem[693] <= 13'b1111111000101;
    mem[694] <= 13'b1101001000010;
    mem[695] <= 13'b1010110101111;
    mem[696] <= 13'b1000111101000;
    mem[697] <= 13'b0111011001000;
    mem[698] <= 13'b0110000110100;
    mem[699] <= 13'b0101000010010;
    mem[700] <= 13'b0100001010001;
    mem[701] <= 13'b0011011011101;
    mem[702] <= 13'b0010110101010;
    mem[703] <= 13'b0010010101100;
    mem[704] <= 13'b0001111011100;
    mem[705] <= 13'b0001100101111;
    mem[706] <= 13'b0001010100001;
    mem[707] <= 13'b0001000101011;
    mem[708] <= 13'b0000111001010;
    mem[709] <= 13'b0000101111010;
    mem[710] <= 13'b0000100111000;
    mem[711] <= 13'b0000100000001;
    mem[712] <= 13'b0000011010100;
    mem[713] <= 13'b0000010101111;
    mem[714] <= 13'b0000010010001;
    mem[715] <= 13'b0000001110111;
    mem[716] <= 13'b0000001100010;
    mem[717] <= 13'b0000001010001;
    mem[718] <= 13'b0000001000011;
    mem[719] <= 13'b0000000110111;
    mem[720] <= 13'b0100000110000;
    mem[721] <= 13'b0001110111100;
    mem[722] <= 13'b0000001100101;
    mem[723] <= 13'b0100100010110;
    mem[724] <= 13'b0010010011100;
    mem[725] <= 13'b1000110110010;
    mem[726] <= 13'b0110011111010;
    mem[727] <= 13'b1011110100110;
    mem[728] <= 13'b1111101111111;
    mem[729] <= 13'b1001010001000;
    mem[730] <= 13'b1101100010101;
    mem[731] <= 13'b0000000000000;
    mem[732] <= 13'b0010011100010;
    mem[733] <= 13'b0101111001001;
    mem[734] <= 13'b1010101111101;
    mem[735] <= 13'b0001000110100;
    mem[736] <= 13'b1000110111001;
    mem[737] <= 13'b0001111010000;
    mem[738] <= 13'b1100000110001;
    mem[739] <= 13'b0111010000110;
    mem[740] <= 13'b0011001110110;
    mem[741] <= 13'b1111111000101;
    mem[742] <= 13'b1101001000010;
    mem[743] <= 13'b1010110101111;
    mem[744] <= 13'b1000111101000;
    mem[745] <= 13'b0111011001000;
    mem[746] <= 13'b0110000110100;
    mem[747] <= 13'b0101000010010;
    mem[748] <= 13'b0100001010001;
    mem[749] <= 13'b0011011011101;
    mem[750] <= 13'b0010110101010;
    mem[751] <= 13'b0010010101100;
    mem[752] <= 13'b0001111011100;
    mem[753] <= 13'b0001100101111;
    mem[754] <= 13'b0001010100001;
    mem[755] <= 13'b0001000101011;
    mem[756] <= 13'b0000111001010;
    mem[757] <= 13'b0000101111010;
    mem[758] <= 13'b0000100111000;
    mem[759] <= 13'b0000100000001;
    mem[760] <= 13'b0000011010100;
    mem[761] <= 13'b0000010101111;
    mem[762] <= 13'b0000010010001;
    mem[763] <= 13'b0000001110111;
    mem[764] <= 13'b0000001100010;
    mem[765] <= 13'b0000001010001;
    mem[766] <= 13'b0000001000011;
    mem[767] <= 13'b0000000110111;
    mem[768] <= 13'b1110101000110;
    mem[769] <= 13'b1000000100010;
    mem[770] <= 13'b0001001100111;
    mem[771] <= 13'b0010111000000;
    mem[772] <= 13'b1010110010011;
    mem[773] <= 13'b1001110111010;
    mem[774] <= 13'b1001100100010;
    mem[775] <= 13'b1111010000111;
    mem[776] <= 13'b1110100000100;
    mem[777] <= 13'b1110100110100;
    mem[778] <= 13'b0110000010111;
    mem[779] <= 13'b1001100001111;
    mem[780] <= 13'b1011110011011;
    mem[781] <= 13'b1110011111101;
    mem[782] <= 13'b0010010110010;
    mem[783] <= 13'b0111101010111;
    mem[784] <= 13'b1110011100100;
    mem[785] <= 13'b0110100110111;
    mem[786] <= 13'b0000000001111;
    mem[787] <= 13'b1010100010100;
    mem[788] <= 13'b0101111101000;
    mem[789] <= 13'b0010001001000;
    mem[790] <= 13'b1110111111110;
    mem[791] <= 13'b1100011000110;
    mem[792] <= 13'b1010001110110;
    mem[793] <= 13'b1000011100100;
    mem[794] <= 13'b0110111110010;
    mem[795] <= 13'b0101110000011;
    mem[796] <= 13'b0100110000001;
    mem[797] <= 13'b0011111011000;
    mem[798] <= 13'b0011001111001;
    mem[799] <= 13'b0010101010111;
    mem[800] <= 13'b0010001101001;
    mem[801] <= 13'b0001110100100;
    mem[802] <= 13'b0001100000001;
    mem[803] <= 13'b0001001111010;
    mem[804] <= 13'b0001000001100;
    mem[805] <= 13'b0000110110000;
    mem[806] <= 13'b0000101100101;
    mem[807] <= 13'b0000100100110;
    mem[808] <= 13'b0000011110011;
    mem[809] <= 13'b0000011001000;
    mem[810] <= 13'b0000010100101;
    mem[811] <= 13'b0000010001000;
    mem[812] <= 13'b0000001110000;
    mem[813] <= 13'b0000001011101;
    mem[814] <= 13'b0000001001100;
    mem[815] <= 13'b0000000111111;
    mem[816] <= 13'b1110101000110;
    mem[817] <= 13'b1000000100010;
    mem[818] <= 13'b0001001100111;
    mem[819] <= 13'b0010111000000;
    mem[820] <= 13'b1010110010011;
    mem[821] <= 13'b1001110111010;
    mem[822] <= 13'b1001100100010;
    mem[823] <= 13'b1111010000111;
    mem[824] <= 13'b1110100000100;
    mem[825] <= 13'b1110100110100;
    mem[826] <= 13'b0110000010111;
    mem[827] <= 13'b1001100001111;
    mem[828] <= 13'b1011110011011;
    mem[829] <= 13'b1110011111101;
    mem[830] <= 13'b0010010110010;
    mem[831] <= 13'b0111101010111;
    mem[832] <= 13'b1110011100100;
    mem[833] <= 13'b0110100110111;
    mem[834] <= 13'b0000000001111;
    mem[835] <= 13'b1010100010100;
    mem[836] <= 13'b0101111101000;
    mem[837] <= 13'b0010001001000;
    mem[838] <= 13'b1110111111110;
    mem[839] <= 13'b1100011000110;
    mem[840] <= 13'b1010001110110;
    mem[841] <= 13'b1000011100100;
    mem[842] <= 13'b0110111110010;
    mem[843] <= 13'b0101110000011;
    mem[844] <= 13'b0100110000001;
    mem[845] <= 13'b0011111011000;
    mem[846] <= 13'b0011001111001;
    mem[847] <= 13'b0010101010111;
    mem[848] <= 13'b0010001101001;
    mem[849] <= 13'b0001110100100;
    mem[850] <= 13'b0001100000001;
    mem[851] <= 13'b0001001111010;
    mem[852] <= 13'b0001000001100;
    mem[853] <= 13'b0000110110000;
    mem[854] <= 13'b0000101100101;
    mem[855] <= 13'b0000100100110;
    mem[856] <= 13'b0000011110011;
    mem[857] <= 13'b0000011001000;
    mem[858] <= 13'b0000010100101;
    mem[859] <= 13'b0000010001000;
    mem[860] <= 13'b0000001110000;
    mem[861] <= 13'b0000001011101;
    mem[862] <= 13'b0000001001100;
    mem[863] <= 13'b0000000111111;
    mem[864] <= 13'b0100110000000;
    mem[865] <= 13'b0100011111101;
    mem[866] <= 13'b1100100001000;
    mem[867] <= 13'b0111110000111;
    mem[868] <= 13'b0001111010010;
    mem[869] <= 13'b1001011100110;
    mem[870] <= 13'b0101010110101;
    mem[871] <= 13'b1011001010110;
    mem[872] <= 13'b0111011010101;
    mem[873] <= 13'b1111111100010;
    mem[874] <= 13'b1100000000110;
    mem[875] <= 13'b0001100000101;
    mem[876] <= 13'b0100001111111;
    mem[877] <= 13'b0110100011111;
    mem[878] <= 13'b1001101001010;
    mem[879] <= 13'b1110000011111;
    mem[880] <= 13'b0011111011100;
    mem[881] <= 13'b1011010000001;
    mem[882] <= 13'b0011111011101;
    mem[883] <= 13'b1101110011001;
    mem[884] <= 13'b1000101010100;
    mem[885] <= 13'b0100011001000;
    mem[886] <= 13'b0000110111000;
    mem[887] <= 13'b1101111011011;
    mem[888] <= 13'b1011100000011;
    mem[889] <= 13'b1001100000000;
    mem[890] <= 13'b0111110101111;
    mem[891] <= 13'b0110011110011;
    mem[892] <= 13'b0101010110001;
    mem[893] <= 13'b0100011010011;
    mem[894] <= 13'b0011101001000;
    mem[895] <= 13'b0011000000010;
    mem[896] <= 13'b0010011110111;
    mem[897] <= 13'b0010000011001;
    mem[898] <= 13'b0001101100001;
    mem[899] <= 13'b0001011001010;
    mem[900] <= 13'b0001001001110;
    mem[901] <= 13'b0000111100110;
    mem[902] <= 13'b0000110010001;
    mem[903] <= 13'b0000101001011;
    mem[904] <= 13'b0000100010001;
    mem[905] <= 13'b0000011100001;
    mem[906] <= 13'b0000010111010;
    mem[907] <= 13'b0000010011001;
    mem[908] <= 13'b0000001111111;
    mem[909] <= 13'b0000001101000;
    mem[910] <= 13'b0000001010110;
    mem[911] <= 13'b0000001000111;
    mem[912] <= 13'b0100110000000;
    mem[913] <= 13'b0100011111101;
    mem[914] <= 13'b1100100001000;
    mem[915] <= 13'b0111110000111;
    mem[916] <= 13'b0001111010010;
    mem[917] <= 13'b1001011100110;
    mem[918] <= 13'b0101010110101;
    mem[919] <= 13'b1011001010110;
    mem[920] <= 13'b0111011010101;
    mem[921] <= 13'b1111111100010;
    mem[922] <= 13'b1100000000110;
    mem[923] <= 13'b0001100000101;
    mem[924] <= 13'b0100001111111;
    mem[925] <= 13'b0110100011111;
    mem[926] <= 13'b1001101001010;
    mem[927] <= 13'b1110000011111;
    mem[928] <= 13'b0011111011100;
    mem[929] <= 13'b1011010000001;
    mem[930] <= 13'b0011111011101;
    mem[931] <= 13'b1101110011001;
    mem[932] <= 13'b1000101010100;
    mem[933] <= 13'b0100011001000;
    mem[934] <= 13'b0000110111000;
    mem[935] <= 13'b1101111011011;
    mem[936] <= 13'b1011100000011;
    mem[937] <= 13'b1001100000000;
    mem[938] <= 13'b0111110101111;
    mem[939] <= 13'b0110011110011;
    mem[940] <= 13'b0101010110001;
    mem[941] <= 13'b0100011010011;
    mem[942] <= 13'b0011101001000;
    mem[943] <= 13'b0011000000010;
    mem[944] <= 13'b0010011110111;
    mem[945] <= 13'b0010000011001;
    mem[946] <= 13'b0001101100001;
    mem[947] <= 13'b0001011001010;
    mem[948] <= 13'b0001001001110;
    mem[949] <= 13'b0000111100110;
    mem[950] <= 13'b0000110010001;
    mem[951] <= 13'b0000101001011;
    mem[952] <= 13'b0000100010001;
    mem[953] <= 13'b0000011100001;
    mem[954] <= 13'b0000010111010;
    mem[955] <= 13'b0000010011001;
    mem[956] <= 13'b0000001111111;
    mem[957] <= 13'b0000001101000;
    mem[958] <= 13'b0000001010110;
    mem[959] <= 13'b0000001000111;
  end


  // Combinational ROM read block
  always@(*)
  begin
    if ( addr >= 1'd0 && addr < 10'd960)
      data_out_t <= mem[addr];
    else
    begin
      data_out_t <= {(13){1'b0}};
    end
  end

  // Output register assignment
  assign data_out = data_out_t;

endmodule



//------> ./rtl_dutmgc_rom_38_64_8_1.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1_2/1117371 Production Release
//  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
// 
//  Generated by:   dr655@ecelinux-16.ece.cornell.edu
//  Generated date: Thu Nov 28 19:53:51 2024
// ----------------------------------------------------------------------

// 
module dutmgc_rom_38_64_8_1 (addr, data_out
);
  input [5:0]addr ;
  output [7:0]data_out ;


  // Constants for ROM dimensions
  parameter n_width    = 8;
  parameter n_size     = 64;
  parameter n_numports = 1;
  parameter n_addr_w   = 6;
  parameter n_inreg    = 0;
  parameter n_outreg   = 0;

  // Declare storage for memory elements
  reg [7:0] mem [63:0];

  // Declare output registers
  reg [7:0] data_out_t;

  // Initialize ROM contents
  initial begin: rom_init_blk
    mem[0] <= 8'b00001010;
    mem[1] <= 8'b00100010;
    mem[2] <= 8'b01100101;
    mem[3] <= 8'b00010010;
    mem[4] <= 8'b00000001;
    mem[5] <= 8'b10101001;
    mem[6] <= 8'b00100001;
    mem[7] <= 8'b01011010;
    mem[8] <= 8'b01010001;
    mem[9] <= 8'b01000101;
    mem[10] <= 8'b00000101;
    mem[11] <= 8'b10010101;
    mem[12] <= 8'b10011010;
    mem[13] <= 8'b10001000;
    mem[14] <= 8'b01011001;
    mem[15] <= 8'b10001001;
    mem[16] <= 8'b10011010;
    mem[17] <= 8'b10101000;
    mem[18] <= 8'b10101010;
    mem[19] <= 8'b01100100;
    mem[20] <= 8'b01001010;
    mem[21] <= 8'b00000101;
    mem[22] <= 8'b01010110;
    mem[23] <= 8'b01010001;
    mem[24] <= 8'b10100110;
    mem[25] <= 8'b00101001;
    mem[26] <= 8'b01000001;
    mem[27] <= 8'b10011001;
    mem[28] <= 8'b00010101;
    mem[29] <= 8'b10101001;
    mem[30] <= 8'b01010110;
    mem[31] <= 8'b10100101;
    mem[32] <= 8'b10101001;
    mem[33] <= 8'b10000010;
    mem[34] <= 8'b00100101;
    mem[35] <= 8'b01010010;
    mem[36] <= 8'b10000010;
    mem[37] <= 8'b01010110;
    mem[38] <= 8'b10010010;
    mem[39] <= 8'b01001000;
    mem[40] <= 8'b10010100;
    mem[41] <= 8'b10010001;
    mem[42] <= 8'b01100101;
    mem[43] <= 8'b01010000;
    mem[44] <= 8'b01011010;
    mem[45] <= 8'b01100001;
    mem[46] <= 8'b01101010;
    mem[47] <= 8'b10100000;
    mem[48] <= 8'b10010000;
    mem[49] <= 8'b01010100;
    mem[50] <= 8'b01010000;
    mem[51] <= 8'b01010101;
    mem[52] <= 8'b01011000;
    mem[53] <= 8'b01001001;
    mem[54] <= 8'b01011001;
    mem[55] <= 8'b00000110;
    mem[56] <= 8'b10000100;
    mem[57] <= 8'b10100110;
    mem[58] <= 8'b10010101;
    mem[59] <= 8'b10000110;
    mem[60] <= 8'b00010110;
    mem[61] <= 8'b10101000;
    mem[62] <= 8'b10100010;
    mem[63] <= 8'b01001010;
  end


  // Combinational ROM read block
  always@(*)
  begin
    data_out_t <= mem[addr];
  end

  // Output register assignment
  assign data_out = data_out_t;

endmodule



//------> ./rtl_dutmgc_rom_39_64_8_1.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1_2/1117371 Production Release
//  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
// 
//  Generated by:   dr655@ecelinux-16.ece.cornell.edu
//  Generated date: Thu Nov 28 19:53:51 2024
// ----------------------------------------------------------------------

// 
module dutmgc_rom_39_64_8_1 (addr, data_out
);
  input [5:0]addr ;
  output [7:0]data_out ;


  // Constants for ROM dimensions
  parameter n_width    = 8;
  parameter n_size     = 64;
  parameter n_numports = 1;
  parameter n_addr_w   = 6;
  parameter n_inreg    = 0;
  parameter n_outreg   = 0;

  // Declare storage for memory elements
  reg [7:0] mem [63:0];

  // Declare output registers
  reg [7:0] data_out_t;

  // Initialize ROM contents
  initial begin: rom_init_blk
    mem[0] <= 8'b10000010;
    mem[1] <= 8'b00011001;
    mem[2] <= 8'b01000101;
    mem[3] <= 8'b10101000;
    mem[4] <= 8'b00011001;
    mem[5] <= 8'b00001010;
    mem[6] <= 8'b10010101;
    mem[7] <= 8'b00010100;
    mem[8] <= 8'b00010101;
    mem[9] <= 8'b10010000;
    mem[10] <= 8'b00001001;
    mem[11] <= 8'b01100010;
    mem[12] <= 8'b10001010;
    mem[13] <= 8'b10010010;
    mem[14] <= 8'b01010001;
    mem[15] <= 8'b01101010;
    mem[16] <= 8'b10100001;
    mem[17] <= 8'b01100110;
    mem[18] <= 8'b00101000;
    mem[19] <= 8'b01010000;
    mem[20] <= 8'b01101000;
    mem[21] <= 8'b00100000;
    mem[22] <= 8'b10100101;
    mem[23] <= 8'b10100100;
    mem[24] <= 8'b10010010;
    mem[25] <= 8'b00000010;
    mem[26] <= 8'b01101000;
    mem[27] <= 8'b10010001;
    mem[28] <= 8'b00101000;
    mem[29] <= 8'b00011010;
    mem[30] <= 8'b10000010;
    mem[31] <= 8'b01011010;
    mem[32] <= 8'b00000010;
    mem[33] <= 8'b00001001;
    mem[34] <= 8'b00000101;
    mem[35] <= 8'b01000101;
    mem[36] <= 8'b10001000;
    mem[37] <= 8'b01100010;
    mem[38] <= 8'b00001001;
    mem[39] <= 8'b10010010;
    mem[40] <= 8'b00000001;
    mem[41] <= 8'b01101001;
    mem[42] <= 8'b01101001;
    mem[43] <= 8'b00100101;
    mem[44] <= 8'b00010100;
    mem[45] <= 8'b00001000;
    mem[46] <= 8'b00101010;
    mem[47] <= 8'b10011010;
    mem[48] <= 8'b00010100;
    mem[49] <= 8'b01101001;
    mem[50] <= 8'b00100110;
    mem[51] <= 8'b10010000;
    mem[52] <= 8'b10001000;
    mem[53] <= 8'b10010000;
    mem[54] <= 8'b00000100;
    mem[55] <= 8'b00010000;
    mem[56] <= 8'b10101000;
    mem[57] <= 8'b00011000;
    mem[58] <= 8'b00000100;
    mem[59] <= 8'b10010000;
    mem[60] <= 8'b01100110;
    mem[61] <= 8'b00011000;
    mem[62] <= 8'b00010000;
    mem[63] <= 8'b00010100;
  end


  // Combinational ROM read block
  always@(*)
  begin
    data_out_t <= mem[addr];
  end

  // Output register assignment
  assign data_out = data_out_t;

endmodule



//------> ./rtl_dutmgc_rom_40_32_19_1.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1_2/1117371 Production Release
//  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
// 
//  Generated by:   dr655@ecelinux-16.ece.cornell.edu
//  Generated date: Thu Nov 28 19:53:51 2024
// ----------------------------------------------------------------------

// 
module dutmgc_rom_40_32_19_1 (addr, data_out
);
  input [4:0]addr ;
  output [18:0]data_out ;


  // Constants for ROM dimensions
  parameter n_width    = 19;
  parameter n_size     = 32;
  parameter n_numports = 1;
  parameter n_addr_w   = 5;
  parameter n_inreg    = 0;
  parameter n_outreg   = 0;

  // Declare storage for memory elements
  reg [18:0] mem [31:0];

  // Declare output registers
  reg [18:0] data_out_t;

  // Initialize ROM contents
  initial begin: rom_init_blk
    mem[0] <= 19'b0000000000101000010;
    mem[1] <= 19'b0000001010001111110;
    mem[2] <= 19'b1111101100100110111;
    mem[3] <= 19'b0000001000110101000;
    mem[4] <= 19'b1111111111101011110;
    mem[5] <= 19'b0000001000001100101;
    mem[6] <= 19'b1111010101010001101;
    mem[7] <= 19'b1111110000100011001;
    mem[8] <= 19'b0000010000001111001;
    mem[9] <= 19'b0000000010101011100;
    mem[10] <= 19'b0000000001111001000;
    mem[11] <= 19'b1111101110010101111;
    mem[12] <= 19'b1010110101101110011;
    mem[13] <= 19'b1111000101010001000;
    mem[14] <= 19'b0011111100000101010;
    mem[15] <= 19'b0010100100101111011;
    mem[16] <= 19'b0000010110011000101;
    mem[17] <= 19'b1111111010101000111;
    mem[18] <= 19'b0000001001001001001;
    mem[19] <= 19'b1111111010011110110;
    mem[20] <= 19'b1100000010011111010;
    mem[21] <= 19'b0010000100001011101;
    mem[22] <= 19'b0010111101010111111;
    mem[23] <= 19'b0100000100000111010;
    mem[24] <= 19'b0000000001100100111;
    mem[25] <= 19'b1111111101111100110;
    mem[26] <= 19'b0000000011011101111;
    mem[27] <= 19'b1111100111111000010;
    mem[28] <= 19'b1110010000011101100;
    mem[29] <= 19'b1110011010101110011;
    mem[30] <= 19'b0011110000011010100;
    mem[31] <= 19'b0001000001000001000;
  end


  // Combinational ROM read block
  always@(*)
  begin
    data_out_t <= mem[addr];
  end

  // Output register assignment
  assign data_out = data_out_t;

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1_2/1117371 Production Release
//  HLS Date:       Fri Jun 28 23:58:31 PDT 2024
// 
//  Generated by:   dr655@ecelinux-16.ece.cornell.edu
//  Generated date: Thu Nov 28 19:53:50 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_16_6_40_48_1_48_40_1_gen
// ------------------------------------------------------------------


module dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_16_6_40_48_1_48_40_1_gen (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [39:0] q;
  output re;
  output [5:0] radr;
  output we;
  output [39:0] d;
  output [5:0] wadr;
  input clken_d;
  input [39:0] d_d;
  output [39:0] q_d;
  input [5:0] radr_d;
  input re_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_15_6_40_48_1_48_40_1_gen
// ------------------------------------------------------------------


module dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_15_6_40_48_1_48_40_1_gen (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [39:0] q;
  output re;
  output [5:0] radr;
  output we;
  output [39:0] d;
  output [5:0] wadr;
  input clken_d;
  input [39:0] d_d;
  output [39:0] q_d;
  input [5:0] radr_d;
  input re_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_14_6_40_48_1_48_40_1_gen
// ------------------------------------------------------------------


module dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_14_6_40_48_1_48_40_1_gen (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [39:0] q;
  output re;
  output [5:0] radr;
  output we;
  output [39:0] d;
  output [5:0] wadr;
  input clken_d;
  input [39:0] d_d;
  output [39:0] q_d;
  input [5:0] radr_d;
  input re_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dut_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module dut_core_core_fsm (
  clk, rst, attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1, fsm_output, for_for_C_2_tr0,
      compute_sqrt_for_C_15_tr0, RMS_NORM_LOOP_2_C_4_tr0, QUANTIZE_ACTIVATION_LOOP_3_C_2_tr0,
      LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0, LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0,
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_63_tr0, RESHAPE_2D_TO_3D_LOOP_3_C_0_tr0, RESHAPE_2D_TO_3D_LOOP_2_C_0_tr0,
      RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0, RESHAPE_2D_TO_3D_LOOP_2_2_C_0_tr0, APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0,
      APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0, CACHE_UPDATE_LOOP_3_C_1_tr0, CACHE_UPDATE_LOOP_2_C_0_tr0,
      CACHE_UPDATE_LOOP_1_C_0_tr0, TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0, TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0,
      TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0, GEMM_3D_FLOAT_LOOP_4_C_3_tr0, GEMM_3D_FLOAT_LOOP_3_C_1_tr0,
      GEMM_3D_FLOAT_LOOP_1_C_0_tr0, SF_LOOP_3_C_0_tr0, SF_LOOP_1_C_0_tr0, CM_LOOP_1_C_0_tr0,
      SOFTMAX_LOOP_3_C_0_tr0, SOFTMAX_LOOP_4_C_2_tr0, SOFTMAX_LOOP_5_C_19_tr0, SOFTMAX_LOOP_1_C_1_tr0,
      GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0, GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0, GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0,
      ATTN_2D_LOOP_3_C_0_tr0, ATTN_2D_LOOP_2_C_0_tr0, RMS_NORM_LOOP_1_2_C_2_tr0,
      compute_sqrt_1_for_C_15_tr0, RMS_NORM_LOOP_2_2_C_4_tr0, QUANTIZE_ACTIVATION_LOOP_3_1_C_2_tr0,
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0, LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0,
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31_tr0, for_1_for_C_1_tr0
);
  input clk;
  input rst;
  input attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1;
  output [8:0] fsm_output;
  reg [8:0] fsm_output;
  input for_for_C_2_tr0;
  input compute_sqrt_for_C_15_tr0;
  input RMS_NORM_LOOP_2_C_4_tr0;
  input QUANTIZE_ACTIVATION_LOOP_3_C_2_tr0;
  input LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0;
  input LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0;
  input LINEAR_FORWARD_NO_MUL_LOOP_2_C_63_tr0;
  input RESHAPE_2D_TO_3D_LOOP_3_C_0_tr0;
  input RESHAPE_2D_TO_3D_LOOP_2_C_0_tr0;
  input RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0;
  input RESHAPE_2D_TO_3D_LOOP_2_2_C_0_tr0;
  input APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0;
  input APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0;
  input CACHE_UPDATE_LOOP_3_C_1_tr0;
  input CACHE_UPDATE_LOOP_2_C_0_tr0;
  input CACHE_UPDATE_LOOP_1_C_0_tr0;
  input TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0;
  input TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0;
  input TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0;
  input GEMM_3D_FLOAT_LOOP_4_C_3_tr0;
  input GEMM_3D_FLOAT_LOOP_3_C_1_tr0;
  input GEMM_3D_FLOAT_LOOP_1_C_0_tr0;
  input SF_LOOP_3_C_0_tr0;
  input SF_LOOP_1_C_0_tr0;
  input CM_LOOP_1_C_0_tr0;
  input SOFTMAX_LOOP_3_C_0_tr0;
  input SOFTMAX_LOOP_4_C_2_tr0;
  input SOFTMAX_LOOP_5_C_19_tr0;
  input SOFTMAX_LOOP_1_C_1_tr0;
  input GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0;
  input GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0;
  input GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0;
  input ATTN_2D_LOOP_3_C_0_tr0;
  input ATTN_2D_LOOP_2_C_0_tr0;
  input RMS_NORM_LOOP_1_2_C_2_tr0;
  input compute_sqrt_1_for_C_15_tr0;
  input RMS_NORM_LOOP_2_2_C_4_tr0;
  input QUANTIZE_ACTIVATION_LOOP_3_1_C_2_tr0;
  input LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0;
  input LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0;
  input LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31_tr0;
  input for_1_for_C_1_tr0;


  // FSM State Type Declaration for dut_core_core_fsm_1
  parameter
    main_C_0 = 9'd0,
    for_for_C_0 = 9'd1,
    for_for_C_1 = 9'd2,
    for_for_C_2 = 9'd3,
    main_C_1 = 9'd4,
    compute_sqrt_for_C_0 = 9'd5,
    compute_sqrt_for_C_1 = 9'd6,
    compute_sqrt_for_C_2 = 9'd7,
    compute_sqrt_for_C_3 = 9'd8,
    compute_sqrt_for_C_4 = 9'd9,
    compute_sqrt_for_C_5 = 9'd10,
    compute_sqrt_for_C_6 = 9'd11,
    compute_sqrt_for_C_7 = 9'd12,
    compute_sqrt_for_C_8 = 9'd13,
    compute_sqrt_for_C_9 = 9'd14,
    compute_sqrt_for_C_10 = 9'd15,
    compute_sqrt_for_C_11 = 9'd16,
    compute_sqrt_for_C_12 = 9'd17,
    compute_sqrt_for_C_13 = 9'd18,
    compute_sqrt_for_C_14 = 9'd19,
    compute_sqrt_for_C_15 = 9'd20,
    main_C_2 = 9'd21,
    main_C_3 = 9'd22,
    main_C_4 = 9'd23,
    main_C_5 = 9'd24,
    main_C_6 = 9'd25,
    main_C_7 = 9'd26,
    main_C_8 = 9'd27,
    main_C_9 = 9'd28,
    main_C_10 = 9'd29,
    main_C_11 = 9'd30,
    main_C_12 = 9'd31,
    main_C_13 = 9'd32,
    main_C_14 = 9'd33,
    main_C_15 = 9'd34,
    main_C_16 = 9'd35,
    main_C_17 = 9'd36,
    main_C_18 = 9'd37,
    main_C_19 = 9'd38,
    main_C_20 = 9'd39,
    main_C_21 = 9'd40,
    main_C_22 = 9'd41,
    main_C_23 = 9'd42,
    main_C_24 = 9'd43,
    main_C_25 = 9'd44,
    main_C_26 = 9'd45,
    main_C_27 = 9'd46,
    main_C_28 = 9'd47,
    main_C_29 = 9'd48,
    main_C_30 = 9'd49,
    main_C_31 = 9'd50,
    main_C_32 = 9'd51,
    main_C_33 = 9'd52,
    RMS_NORM_LOOP_2_C_0 = 9'd53,
    RMS_NORM_LOOP_2_C_1 = 9'd54,
    RMS_NORM_LOOP_2_C_2 = 9'd55,
    RMS_NORM_LOOP_2_C_3 = 9'd56,
    RMS_NORM_LOOP_2_C_4 = 9'd57,
    main_C_34 = 9'd58,
    main_C_35 = 9'd59,
    main_C_36 = 9'd60,
    main_C_37 = 9'd61,
    main_C_38 = 9'd62,
    main_C_39 = 9'd63,
    main_C_40 = 9'd64,
    main_C_41 = 9'd65,
    main_C_42 = 9'd66,
    main_C_43 = 9'd67,
    main_C_44 = 9'd68,
    main_C_45 = 9'd69,
    main_C_46 = 9'd70,
    main_C_47 = 9'd71,
    main_C_48 = 9'd72,
    QUANTIZE_ACTIVATION_LOOP_3_C_0 = 9'd73,
    QUANTIZE_ACTIVATION_LOOP_3_C_1 = 9'd74,
    QUANTIZE_ACTIVATION_LOOP_3_C_2 = 9'd75,
    LINEAR_FORWARD_NO_MUL_LOOP_3_C_0 = 9'd76,
    LINEAR_FORWARD_NO_MUL_LOOP_4_C_0 = 9'd77,
    LINEAR_FORWARD_NO_MUL_LOOP_3_C_1 = 9'd78,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_0 = 9'd79,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_1 = 9'd80,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_2 = 9'd81,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_3 = 9'd82,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_4 = 9'd83,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_5 = 9'd84,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_6 = 9'd85,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_7 = 9'd86,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_8 = 9'd87,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_9 = 9'd88,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_10 = 9'd89,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_11 = 9'd90,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_12 = 9'd91,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_13 = 9'd92,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_14 = 9'd93,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_15 = 9'd94,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_16 = 9'd95,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_17 = 9'd96,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_18 = 9'd97,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_19 = 9'd98,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_20 = 9'd99,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_21 = 9'd100,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_22 = 9'd101,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_23 = 9'd102,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_24 = 9'd103,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_25 = 9'd104,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_26 = 9'd105,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_27 = 9'd106,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_28 = 9'd107,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_29 = 9'd108,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_30 = 9'd109,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_31 = 9'd110,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_32 = 9'd111,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_33 = 9'd112,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_34 = 9'd113,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_35 = 9'd114,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_36 = 9'd115,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_37 = 9'd116,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_38 = 9'd117,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_39 = 9'd118,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_40 = 9'd119,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_41 = 9'd120,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_42 = 9'd121,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_43 = 9'd122,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_44 = 9'd123,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_45 = 9'd124,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_46 = 9'd125,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_47 = 9'd126,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_48 = 9'd127,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_49 = 9'd128,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_50 = 9'd129,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_51 = 9'd130,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_52 = 9'd131,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_53 = 9'd132,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_54 = 9'd133,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_55 = 9'd134,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_56 = 9'd135,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_57 = 9'd136,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_58 = 9'd137,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_59 = 9'd138,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_60 = 9'd139,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_61 = 9'd140,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_62 = 9'd141,
    LINEAR_FORWARD_NO_MUL_LOOP_2_C_63 = 9'd142,
    RESHAPE_2D_TO_3D_LOOP_3_C_0 = 9'd143,
    RESHAPE_2D_TO_3D_LOOP_2_C_0 = 9'd144,
    RESHAPE_2D_TO_3D_LOOP_3_2_C_0 = 9'd145,
    RESHAPE_2D_TO_3D_LOOP_2_2_C_0 = 9'd146,
    APPLY_ROTARY_POS_EMB_LOOP_6_C_0 = 9'd147,
    APPLY_ROTARY_POS_EMB_LOOP_6_C_1 = 9'd148,
    APPLY_ROTARY_POS_EMB_LOOP_6_C_2 = 9'd149,
    APPLY_ROTARY_POS_EMB_LOOP_4_C_0 = 9'd150,
    CACHE_UPDATE_LOOP_3_C_0 = 9'd151,
    CACHE_UPDATE_LOOP_3_C_1 = 9'd152,
    CACHE_UPDATE_LOOP_2_C_0 = 9'd153,
    CACHE_UPDATE_LOOP_1_C_0 = 9'd154,
    TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_0 = 9'd155,
    TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_1 = 9'd156,
    TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2 = 9'd157,
    TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0 = 9'd158,
    TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0 = 9'd159,
    GEMM_3D_FLOAT_LOOP_3_C_0 = 9'd160,
    GEMM_3D_FLOAT_LOOP_4_C_0 = 9'd161,
    GEMM_3D_FLOAT_LOOP_4_C_1 = 9'd162,
    GEMM_3D_FLOAT_LOOP_4_C_2 = 9'd163,
    GEMM_3D_FLOAT_LOOP_4_C_3 = 9'd164,
    GEMM_3D_FLOAT_LOOP_3_C_1 = 9'd165,
    GEMM_3D_FLOAT_LOOP_1_C_0 = 9'd166,
    SF_LOOP_3_C_0 = 9'd167,
    SF_LOOP_1_C_0 = 9'd168,
    CM_LOOP_1_C_0 = 9'd169,
    SOFTMAX_LOOP_1_C_0 = 9'd170,
    SOFTMAX_LOOP_3_C_0 = 9'd171,
    SOFTMAX_LOOP_4_C_0 = 9'd172,
    SOFTMAX_LOOP_4_C_1 = 9'd173,
    SOFTMAX_LOOP_4_C_2 = 9'd174,
    SOFTMAX_LOOP_5_C_0 = 9'd175,
    SOFTMAX_LOOP_5_C_1 = 9'd176,
    SOFTMAX_LOOP_5_C_2 = 9'd177,
    SOFTMAX_LOOP_5_C_3 = 9'd178,
    SOFTMAX_LOOP_5_C_4 = 9'd179,
    SOFTMAX_LOOP_5_C_5 = 9'd180,
    SOFTMAX_LOOP_5_C_6 = 9'd181,
    SOFTMAX_LOOP_5_C_7 = 9'd182,
    SOFTMAX_LOOP_5_C_8 = 9'd183,
    SOFTMAX_LOOP_5_C_9 = 9'd184,
    SOFTMAX_LOOP_5_C_10 = 9'd185,
    SOFTMAX_LOOP_5_C_11 = 9'd186,
    SOFTMAX_LOOP_5_C_12 = 9'd187,
    SOFTMAX_LOOP_5_C_13 = 9'd188,
    SOFTMAX_LOOP_5_C_14 = 9'd189,
    SOFTMAX_LOOP_5_C_15 = 9'd190,
    SOFTMAX_LOOP_5_C_16 = 9'd191,
    SOFTMAX_LOOP_5_C_17 = 9'd192,
    SOFTMAX_LOOP_5_C_18 = 9'd193,
    SOFTMAX_LOOP_5_C_19 = 9'd194,
    SOFTMAX_LOOP_1_C_1 = 9'd195,
    GEMM_3D_FLOAT_LOOP_3_1_C_0 = 9'd196,
    GEMM_3D_FLOAT_LOOP_4_1_C_0 = 9'd197,
    GEMM_3D_FLOAT_LOOP_4_1_C_1 = 9'd198,
    GEMM_3D_FLOAT_LOOP_4_1_C_2 = 9'd199,
    GEMM_3D_FLOAT_LOOP_4_1_C_3 = 9'd200,
    GEMM_3D_FLOAT_LOOP_3_1_C_1 = 9'd201,
    GEMM_3D_FLOAT_LOOP_1_1_C_0 = 9'd202,
    ATTN_2D_LOOP_3_C_0 = 9'd203,
    ATTN_2D_LOOP_2_C_0 = 9'd204,
    RMS_NORM_LOOP_1_2_C_0 = 9'd205,
    RMS_NORM_LOOP_1_2_C_1 = 9'd206,
    RMS_NORM_LOOP_1_2_C_2 = 9'd207,
    main_C_49 = 9'd208,
    compute_sqrt_1_for_C_0 = 9'd209,
    compute_sqrt_1_for_C_1 = 9'd210,
    compute_sqrt_1_for_C_2 = 9'd211,
    compute_sqrt_1_for_C_3 = 9'd212,
    compute_sqrt_1_for_C_4 = 9'd213,
    compute_sqrt_1_for_C_5 = 9'd214,
    compute_sqrt_1_for_C_6 = 9'd215,
    compute_sqrt_1_for_C_7 = 9'd216,
    compute_sqrt_1_for_C_8 = 9'd217,
    compute_sqrt_1_for_C_9 = 9'd218,
    compute_sqrt_1_for_C_10 = 9'd219,
    compute_sqrt_1_for_C_11 = 9'd220,
    compute_sqrt_1_for_C_12 = 9'd221,
    compute_sqrt_1_for_C_13 = 9'd222,
    compute_sqrt_1_for_C_14 = 9'd223,
    compute_sqrt_1_for_C_15 = 9'd224,
    main_C_50 = 9'd225,
    main_C_51 = 9'd226,
    main_C_52 = 9'd227,
    main_C_53 = 9'd228,
    main_C_54 = 9'd229,
    main_C_55 = 9'd230,
    main_C_56 = 9'd231,
    main_C_57 = 9'd232,
    main_C_58 = 9'd233,
    main_C_59 = 9'd234,
    main_C_60 = 9'd235,
    main_C_61 = 9'd236,
    main_C_62 = 9'd237,
    main_C_63 = 9'd238,
    main_C_64 = 9'd239,
    main_C_65 = 9'd240,
    main_C_66 = 9'd241,
    main_C_67 = 9'd242,
    main_C_68 = 9'd243,
    RMS_NORM_LOOP_2_2_C_0 = 9'd244,
    RMS_NORM_LOOP_2_2_C_1 = 9'd245,
    RMS_NORM_LOOP_2_2_C_2 = 9'd246,
    RMS_NORM_LOOP_2_2_C_3 = 9'd247,
    RMS_NORM_LOOP_2_2_C_4 = 9'd248,
    main_C_69 = 9'd249,
    main_C_70 = 9'd250,
    main_C_71 = 9'd251,
    main_C_72 = 9'd252,
    main_C_73 = 9'd253,
    main_C_74 = 9'd254,
    main_C_75 = 9'd255,
    main_C_76 = 9'd256,
    main_C_77 = 9'd257,
    main_C_78 = 9'd258,
    main_C_79 = 9'd259,
    main_C_80 = 9'd260,
    main_C_81 = 9'd261,
    main_C_82 = 9'd262,
    main_C_83 = 9'd263,
    main_C_84 = 9'd264,
    main_C_85 = 9'd265,
    main_C_86 = 9'd266,
    main_C_87 = 9'd267,
    main_C_88 = 9'd268,
    main_C_89 = 9'd269,
    main_C_90 = 9'd270,
    main_C_91 = 9'd271,
    main_C_92 = 9'd272,
    main_C_93 = 9'd273,
    main_C_94 = 9'd274,
    main_C_95 = 9'd275,
    main_C_96 = 9'd276,
    main_C_97 = 9'd277,
    main_C_98 = 9'd278,
    main_C_99 = 9'd279,
    main_C_100 = 9'd280,
    QUANTIZE_ACTIVATION_LOOP_3_1_C_0 = 9'd281,
    QUANTIZE_ACTIVATION_LOOP_3_1_C_1 = 9'd282,
    QUANTIZE_ACTIVATION_LOOP_3_1_C_2 = 9'd283,
    LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_0 = 9'd284,
    LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0 = 9'd285,
    LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1 = 9'd286,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_0 = 9'd287,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_1 = 9'd288,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_2 = 9'd289,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_3 = 9'd290,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_4 = 9'd291,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_5 = 9'd292,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_6 = 9'd293,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_7 = 9'd294,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_8 = 9'd295,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_9 = 9'd296,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_10 = 9'd297,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_11 = 9'd298,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_12 = 9'd299,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_13 = 9'd300,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_14 = 9'd301,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_15 = 9'd302,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_16 = 9'd303,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_17 = 9'd304,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_18 = 9'd305,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_19 = 9'd306,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_20 = 9'd307,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_21 = 9'd308,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_22 = 9'd309,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_23 = 9'd310,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_24 = 9'd311,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_25 = 9'd312,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_26 = 9'd313,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_27 = 9'd314,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_28 = 9'd315,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_29 = 9'd316,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_30 = 9'd317,
    LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31 = 9'd318,
    for_1_for_C_0 = 9'd319,
    for_1_for_C_1 = 9'd320;

  reg [8:0] state_var;
  reg [8:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : dut_core_core_fsm_1
    case (state_var)
      for_for_C_0 : begin
        fsm_output = 9'b000000001;
        state_var_NS = for_for_C_1;
      end
      for_for_C_1 : begin
        fsm_output = 9'b000000010;
        state_var_NS = for_for_C_2;
      end
      for_for_C_2 : begin
        fsm_output = 9'b000000011;
        if ( for_for_C_2_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_for_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 9'b000000100;
        state_var_NS = compute_sqrt_for_C_0;
      end
      compute_sqrt_for_C_0 : begin
        fsm_output = 9'b000000101;
        state_var_NS = compute_sqrt_for_C_1;
      end
      compute_sqrt_for_C_1 : begin
        fsm_output = 9'b000000110;
        state_var_NS = compute_sqrt_for_C_2;
      end
      compute_sqrt_for_C_2 : begin
        fsm_output = 9'b000000111;
        state_var_NS = compute_sqrt_for_C_3;
      end
      compute_sqrt_for_C_3 : begin
        fsm_output = 9'b000001000;
        state_var_NS = compute_sqrt_for_C_4;
      end
      compute_sqrt_for_C_4 : begin
        fsm_output = 9'b000001001;
        state_var_NS = compute_sqrt_for_C_5;
      end
      compute_sqrt_for_C_5 : begin
        fsm_output = 9'b000001010;
        state_var_NS = compute_sqrt_for_C_6;
      end
      compute_sqrt_for_C_6 : begin
        fsm_output = 9'b000001011;
        state_var_NS = compute_sqrt_for_C_7;
      end
      compute_sqrt_for_C_7 : begin
        fsm_output = 9'b000001100;
        state_var_NS = compute_sqrt_for_C_8;
      end
      compute_sqrt_for_C_8 : begin
        fsm_output = 9'b000001101;
        state_var_NS = compute_sqrt_for_C_9;
      end
      compute_sqrt_for_C_9 : begin
        fsm_output = 9'b000001110;
        state_var_NS = compute_sqrt_for_C_10;
      end
      compute_sqrt_for_C_10 : begin
        fsm_output = 9'b000001111;
        state_var_NS = compute_sqrt_for_C_11;
      end
      compute_sqrt_for_C_11 : begin
        fsm_output = 9'b000010000;
        state_var_NS = compute_sqrt_for_C_12;
      end
      compute_sqrt_for_C_12 : begin
        fsm_output = 9'b000010001;
        state_var_NS = compute_sqrt_for_C_13;
      end
      compute_sqrt_for_C_13 : begin
        fsm_output = 9'b000010010;
        state_var_NS = compute_sqrt_for_C_14;
      end
      compute_sqrt_for_C_14 : begin
        fsm_output = 9'b000010011;
        state_var_NS = compute_sqrt_for_C_15;
      end
      compute_sqrt_for_C_15 : begin
        fsm_output = 9'b000010100;
        if ( compute_sqrt_for_C_15_tr0 ) begin
          state_var_NS = main_C_2;
        end
        else begin
          state_var_NS = compute_sqrt_for_C_0;
        end
      end
      main_C_2 : begin
        fsm_output = 9'b000010101;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 9'b000010110;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 9'b000010111;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 9'b000011000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 9'b000011001;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 9'b000011010;
        state_var_NS = main_C_8;
      end
      main_C_8 : begin
        fsm_output = 9'b000011011;
        state_var_NS = main_C_9;
      end
      main_C_9 : begin
        fsm_output = 9'b000011100;
        state_var_NS = main_C_10;
      end
      main_C_10 : begin
        fsm_output = 9'b000011101;
        state_var_NS = main_C_11;
      end
      main_C_11 : begin
        fsm_output = 9'b000011110;
        state_var_NS = main_C_12;
      end
      main_C_12 : begin
        fsm_output = 9'b000011111;
        state_var_NS = main_C_13;
      end
      main_C_13 : begin
        fsm_output = 9'b000100000;
        state_var_NS = main_C_14;
      end
      main_C_14 : begin
        fsm_output = 9'b000100001;
        state_var_NS = main_C_15;
      end
      main_C_15 : begin
        fsm_output = 9'b000100010;
        state_var_NS = main_C_16;
      end
      main_C_16 : begin
        fsm_output = 9'b000100011;
        state_var_NS = main_C_17;
      end
      main_C_17 : begin
        fsm_output = 9'b000100100;
        state_var_NS = main_C_18;
      end
      main_C_18 : begin
        fsm_output = 9'b000100101;
        state_var_NS = main_C_19;
      end
      main_C_19 : begin
        fsm_output = 9'b000100110;
        state_var_NS = main_C_20;
      end
      main_C_20 : begin
        fsm_output = 9'b000100111;
        state_var_NS = main_C_21;
      end
      main_C_21 : begin
        fsm_output = 9'b000101000;
        state_var_NS = main_C_22;
      end
      main_C_22 : begin
        fsm_output = 9'b000101001;
        state_var_NS = main_C_23;
      end
      main_C_23 : begin
        fsm_output = 9'b000101010;
        state_var_NS = main_C_24;
      end
      main_C_24 : begin
        fsm_output = 9'b000101011;
        state_var_NS = main_C_25;
      end
      main_C_25 : begin
        fsm_output = 9'b000101100;
        state_var_NS = main_C_26;
      end
      main_C_26 : begin
        fsm_output = 9'b000101101;
        state_var_NS = main_C_27;
      end
      main_C_27 : begin
        fsm_output = 9'b000101110;
        state_var_NS = main_C_28;
      end
      main_C_28 : begin
        fsm_output = 9'b000101111;
        state_var_NS = main_C_29;
      end
      main_C_29 : begin
        fsm_output = 9'b000110000;
        state_var_NS = main_C_30;
      end
      main_C_30 : begin
        fsm_output = 9'b000110001;
        state_var_NS = main_C_31;
      end
      main_C_31 : begin
        fsm_output = 9'b000110010;
        state_var_NS = main_C_32;
      end
      main_C_32 : begin
        fsm_output = 9'b000110011;
        state_var_NS = main_C_33;
      end
      main_C_33 : begin
        fsm_output = 9'b000110100;
        state_var_NS = RMS_NORM_LOOP_2_C_0;
      end
      RMS_NORM_LOOP_2_C_0 : begin
        fsm_output = 9'b000110101;
        state_var_NS = RMS_NORM_LOOP_2_C_1;
      end
      RMS_NORM_LOOP_2_C_1 : begin
        fsm_output = 9'b000110110;
        state_var_NS = RMS_NORM_LOOP_2_C_2;
      end
      RMS_NORM_LOOP_2_C_2 : begin
        fsm_output = 9'b000110111;
        state_var_NS = RMS_NORM_LOOP_2_C_3;
      end
      RMS_NORM_LOOP_2_C_3 : begin
        fsm_output = 9'b000111000;
        state_var_NS = RMS_NORM_LOOP_2_C_4;
      end
      RMS_NORM_LOOP_2_C_4 : begin
        fsm_output = 9'b000111001;
        if ( RMS_NORM_LOOP_2_C_4_tr0 ) begin
          state_var_NS = main_C_34;
        end
        else begin
          state_var_NS = RMS_NORM_LOOP_2_C_0;
        end
      end
      main_C_34 : begin
        fsm_output = 9'b000111010;
        state_var_NS = main_C_35;
      end
      main_C_35 : begin
        fsm_output = 9'b000111011;
        state_var_NS = main_C_36;
      end
      main_C_36 : begin
        fsm_output = 9'b000111100;
        state_var_NS = main_C_37;
      end
      main_C_37 : begin
        fsm_output = 9'b000111101;
        state_var_NS = main_C_38;
      end
      main_C_38 : begin
        fsm_output = 9'b000111110;
        state_var_NS = main_C_39;
      end
      main_C_39 : begin
        fsm_output = 9'b000111111;
        state_var_NS = main_C_40;
      end
      main_C_40 : begin
        fsm_output = 9'b001000000;
        state_var_NS = main_C_41;
      end
      main_C_41 : begin
        fsm_output = 9'b001000001;
        state_var_NS = main_C_42;
      end
      main_C_42 : begin
        fsm_output = 9'b001000010;
        state_var_NS = main_C_43;
      end
      main_C_43 : begin
        fsm_output = 9'b001000011;
        state_var_NS = main_C_44;
      end
      main_C_44 : begin
        fsm_output = 9'b001000100;
        state_var_NS = main_C_45;
      end
      main_C_45 : begin
        fsm_output = 9'b001000101;
        state_var_NS = main_C_46;
      end
      main_C_46 : begin
        fsm_output = 9'b001000110;
        state_var_NS = main_C_47;
      end
      main_C_47 : begin
        fsm_output = 9'b001000111;
        state_var_NS = main_C_48;
      end
      main_C_48 : begin
        fsm_output = 9'b001001000;
        state_var_NS = QUANTIZE_ACTIVATION_LOOP_3_C_0;
      end
      QUANTIZE_ACTIVATION_LOOP_3_C_0 : begin
        fsm_output = 9'b001001001;
        state_var_NS = QUANTIZE_ACTIVATION_LOOP_3_C_1;
      end
      QUANTIZE_ACTIVATION_LOOP_3_C_1 : begin
        fsm_output = 9'b001001010;
        state_var_NS = QUANTIZE_ACTIVATION_LOOP_3_C_2;
      end
      QUANTIZE_ACTIVATION_LOOP_3_C_2 : begin
        fsm_output = 9'b001001011;
        if ( QUANTIZE_ACTIVATION_LOOP_3_C_2_tr0 ) begin
          state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_3_C_0;
        end
        else begin
          state_var_NS = QUANTIZE_ACTIVATION_LOOP_3_C_0;
        end
      end
      LINEAR_FORWARD_NO_MUL_LOOP_3_C_0 : begin
        fsm_output = 9'b001001100;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_4_C_0;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_4_C_0 : begin
        fsm_output = 9'b001001101;
        if ( LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0 ) begin
          state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_3_C_1;
        end
        else begin
          state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_4_C_0;
        end
      end
      LINEAR_FORWARD_NO_MUL_LOOP_3_C_1 : begin
        fsm_output = 9'b001001110;
        if ( LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0 ) begin
          state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_0;
        end
        else begin
          state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_3_C_0;
        end
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_0 : begin
        fsm_output = 9'b001001111;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_1;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_1 : begin
        fsm_output = 9'b001010000;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_2;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_2 : begin
        fsm_output = 9'b001010001;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_3;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_3 : begin
        fsm_output = 9'b001010010;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_4;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_4 : begin
        fsm_output = 9'b001010011;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_5;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_5 : begin
        fsm_output = 9'b001010100;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_6;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_6 : begin
        fsm_output = 9'b001010101;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_7;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_7 : begin
        fsm_output = 9'b001010110;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_8;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_8 : begin
        fsm_output = 9'b001010111;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_9;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_9 : begin
        fsm_output = 9'b001011000;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_10;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_10 : begin
        fsm_output = 9'b001011001;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_11;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_11 : begin
        fsm_output = 9'b001011010;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_12;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_12 : begin
        fsm_output = 9'b001011011;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_13;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_13 : begin
        fsm_output = 9'b001011100;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_14;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_14 : begin
        fsm_output = 9'b001011101;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_15;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_15 : begin
        fsm_output = 9'b001011110;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_16;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_16 : begin
        fsm_output = 9'b001011111;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_17;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_17 : begin
        fsm_output = 9'b001100000;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_18;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_18 : begin
        fsm_output = 9'b001100001;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_19;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_19 : begin
        fsm_output = 9'b001100010;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_20;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_20 : begin
        fsm_output = 9'b001100011;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_21;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_21 : begin
        fsm_output = 9'b001100100;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_22;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_22 : begin
        fsm_output = 9'b001100101;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_23;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_23 : begin
        fsm_output = 9'b001100110;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_24;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_24 : begin
        fsm_output = 9'b001100111;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_25;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_25 : begin
        fsm_output = 9'b001101000;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_26;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_26 : begin
        fsm_output = 9'b001101001;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_27;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_27 : begin
        fsm_output = 9'b001101010;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_28;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_28 : begin
        fsm_output = 9'b001101011;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_29;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_29 : begin
        fsm_output = 9'b001101100;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_30;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_30 : begin
        fsm_output = 9'b001101101;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_31;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_31 : begin
        fsm_output = 9'b001101110;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_32;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_32 : begin
        fsm_output = 9'b001101111;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_33;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_33 : begin
        fsm_output = 9'b001110000;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_34;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_34 : begin
        fsm_output = 9'b001110001;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_35;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_35 : begin
        fsm_output = 9'b001110010;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_36;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_36 : begin
        fsm_output = 9'b001110011;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_37;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_37 : begin
        fsm_output = 9'b001110100;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_38;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_38 : begin
        fsm_output = 9'b001110101;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_39;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_39 : begin
        fsm_output = 9'b001110110;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_40;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_40 : begin
        fsm_output = 9'b001110111;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_41;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_41 : begin
        fsm_output = 9'b001111000;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_42;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_42 : begin
        fsm_output = 9'b001111001;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_43;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_43 : begin
        fsm_output = 9'b001111010;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_44;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_44 : begin
        fsm_output = 9'b001111011;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_45;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_45 : begin
        fsm_output = 9'b001111100;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_46;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_46 : begin
        fsm_output = 9'b001111101;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_47;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_47 : begin
        fsm_output = 9'b001111110;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_48;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_48 : begin
        fsm_output = 9'b001111111;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_49;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_49 : begin
        fsm_output = 9'b010000000;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_50;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_50 : begin
        fsm_output = 9'b010000001;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_51;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_51 : begin
        fsm_output = 9'b010000010;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_52;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_52 : begin
        fsm_output = 9'b010000011;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_53;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_53 : begin
        fsm_output = 9'b010000100;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_54;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_54 : begin
        fsm_output = 9'b010000101;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_55;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_55 : begin
        fsm_output = 9'b010000110;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_56;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_56 : begin
        fsm_output = 9'b010000111;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_57;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_57 : begin
        fsm_output = 9'b010001000;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_58;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_58 : begin
        fsm_output = 9'b010001001;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_59;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_59 : begin
        fsm_output = 9'b010001010;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_60;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_60 : begin
        fsm_output = 9'b010001011;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_61;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_61 : begin
        fsm_output = 9'b010001100;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_62;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_62 : begin
        fsm_output = 9'b010001101;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_C_63;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_C_63 : begin
        fsm_output = 9'b010001110;
        if ( LINEAR_FORWARD_NO_MUL_LOOP_2_C_63_tr0 ) begin
          state_var_NS = RESHAPE_2D_TO_3D_LOOP_3_C_0;
        end
        else begin
          state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_3_C_0;
        end
      end
      RESHAPE_2D_TO_3D_LOOP_3_C_0 : begin
        fsm_output = 9'b010001111;
        if ( RESHAPE_2D_TO_3D_LOOP_3_C_0_tr0 ) begin
          state_var_NS = RESHAPE_2D_TO_3D_LOOP_2_C_0;
        end
        else begin
          state_var_NS = RESHAPE_2D_TO_3D_LOOP_3_C_0;
        end
      end
      RESHAPE_2D_TO_3D_LOOP_2_C_0 : begin
        fsm_output = 9'b010010000;
        if ( RESHAPE_2D_TO_3D_LOOP_2_C_0_tr0 ) begin
          state_var_NS = RESHAPE_2D_TO_3D_LOOP_3_2_C_0;
        end
        else begin
          state_var_NS = RESHAPE_2D_TO_3D_LOOP_3_C_0;
        end
      end
      RESHAPE_2D_TO_3D_LOOP_3_2_C_0 : begin
        fsm_output = 9'b010010001;
        if ( RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0 ) begin
          state_var_NS = RESHAPE_2D_TO_3D_LOOP_2_2_C_0;
        end
        else begin
          state_var_NS = RESHAPE_2D_TO_3D_LOOP_3_2_C_0;
        end
      end
      RESHAPE_2D_TO_3D_LOOP_2_2_C_0 : begin
        fsm_output = 9'b010010010;
        if ( RESHAPE_2D_TO_3D_LOOP_2_2_C_0_tr0 ) begin
          state_var_NS = APPLY_ROTARY_POS_EMB_LOOP_6_C_0;
        end
        else begin
          state_var_NS = RESHAPE_2D_TO_3D_LOOP_3_2_C_0;
        end
      end
      APPLY_ROTARY_POS_EMB_LOOP_6_C_0 : begin
        fsm_output = 9'b010010011;
        state_var_NS = APPLY_ROTARY_POS_EMB_LOOP_6_C_1;
      end
      APPLY_ROTARY_POS_EMB_LOOP_6_C_1 : begin
        fsm_output = 9'b010010100;
        state_var_NS = APPLY_ROTARY_POS_EMB_LOOP_6_C_2;
      end
      APPLY_ROTARY_POS_EMB_LOOP_6_C_2 : begin
        fsm_output = 9'b010010101;
        if ( APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0 ) begin
          state_var_NS = APPLY_ROTARY_POS_EMB_LOOP_4_C_0;
        end
        else begin
          state_var_NS = APPLY_ROTARY_POS_EMB_LOOP_6_C_0;
        end
      end
      APPLY_ROTARY_POS_EMB_LOOP_4_C_0 : begin
        fsm_output = 9'b010010110;
        if ( APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0 ) begin
          state_var_NS = CACHE_UPDATE_LOOP_3_C_0;
        end
        else begin
          state_var_NS = APPLY_ROTARY_POS_EMB_LOOP_6_C_0;
        end
      end
      CACHE_UPDATE_LOOP_3_C_0 : begin
        fsm_output = 9'b010010111;
        state_var_NS = CACHE_UPDATE_LOOP_3_C_1;
      end
      CACHE_UPDATE_LOOP_3_C_1 : begin
        fsm_output = 9'b010011000;
        if ( CACHE_UPDATE_LOOP_3_C_1_tr0 ) begin
          state_var_NS = CACHE_UPDATE_LOOP_2_C_0;
        end
        else begin
          state_var_NS = CACHE_UPDATE_LOOP_3_C_0;
        end
      end
      CACHE_UPDATE_LOOP_2_C_0 : begin
        fsm_output = 9'b010011001;
        if ( CACHE_UPDATE_LOOP_2_C_0_tr0 ) begin
          state_var_NS = CACHE_UPDATE_LOOP_1_C_0;
        end
        else begin
          state_var_NS = CACHE_UPDATE_LOOP_3_C_0;
        end
      end
      CACHE_UPDATE_LOOP_1_C_0 : begin
        fsm_output = 9'b010011010;
        if ( CACHE_UPDATE_LOOP_1_C_0_tr0 ) begin
          state_var_NS = TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_0;
        end
        else begin
          state_var_NS = CACHE_UPDATE_LOOP_3_C_0;
        end
      end
      TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_0 : begin
        fsm_output = 9'b010011011;
        state_var_NS = TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_1;
      end
      TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_1 : begin
        fsm_output = 9'b010011100;
        state_var_NS = TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2;
      end
      TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2 : begin
        fsm_output = 9'b010011101;
        if ( TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0 ) begin
          state_var_NS = TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0;
        end
        else begin
          state_var_NS = TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_0;
        end
      end
      TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0 : begin
        fsm_output = 9'b010011110;
        if ( TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0 ) begin
          state_var_NS = TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0;
        end
        else begin
          state_var_NS = TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_0;
        end
      end
      TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0 : begin
        fsm_output = 9'b010011111;
        if ( TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0 ) begin
          state_var_NS = GEMM_3D_FLOAT_LOOP_3_C_0;
        end
        else begin
          state_var_NS = TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_0;
        end
      end
      GEMM_3D_FLOAT_LOOP_3_C_0 : begin
        fsm_output = 9'b010100000;
        state_var_NS = GEMM_3D_FLOAT_LOOP_4_C_0;
      end
      GEMM_3D_FLOAT_LOOP_4_C_0 : begin
        fsm_output = 9'b010100001;
        state_var_NS = GEMM_3D_FLOAT_LOOP_4_C_1;
      end
      GEMM_3D_FLOAT_LOOP_4_C_1 : begin
        fsm_output = 9'b010100010;
        state_var_NS = GEMM_3D_FLOAT_LOOP_4_C_2;
      end
      GEMM_3D_FLOAT_LOOP_4_C_2 : begin
        fsm_output = 9'b010100011;
        state_var_NS = GEMM_3D_FLOAT_LOOP_4_C_3;
      end
      GEMM_3D_FLOAT_LOOP_4_C_3 : begin
        fsm_output = 9'b010100100;
        if ( GEMM_3D_FLOAT_LOOP_4_C_3_tr0 ) begin
          state_var_NS = GEMM_3D_FLOAT_LOOP_3_C_1;
        end
        else begin
          state_var_NS = GEMM_3D_FLOAT_LOOP_4_C_0;
        end
      end
      GEMM_3D_FLOAT_LOOP_3_C_1 : begin
        fsm_output = 9'b010100101;
        if ( GEMM_3D_FLOAT_LOOP_3_C_1_tr0 ) begin
          state_var_NS = GEMM_3D_FLOAT_LOOP_1_C_0;
        end
        else begin
          state_var_NS = GEMM_3D_FLOAT_LOOP_3_C_0;
        end
      end
      GEMM_3D_FLOAT_LOOP_1_C_0 : begin
        fsm_output = 9'b010100110;
        if ( GEMM_3D_FLOAT_LOOP_1_C_0_tr0 ) begin
          state_var_NS = SF_LOOP_3_C_0;
        end
        else begin
          state_var_NS = GEMM_3D_FLOAT_LOOP_3_C_0;
        end
      end
      SF_LOOP_3_C_0 : begin
        fsm_output = 9'b010100111;
        if ( SF_LOOP_3_C_0_tr0 ) begin
          state_var_NS = SF_LOOP_1_C_0;
        end
        else begin
          state_var_NS = SF_LOOP_3_C_0;
        end
      end
      SF_LOOP_1_C_0 : begin
        fsm_output = 9'b010101000;
        if ( SF_LOOP_1_C_0_tr0 ) begin
          state_var_NS = CM_LOOP_1_C_0;
        end
        else begin
          state_var_NS = SF_LOOP_3_C_0;
        end
      end
      CM_LOOP_1_C_0 : begin
        fsm_output = 9'b010101001;
        if ( CM_LOOP_1_C_0_tr0 ) begin
          state_var_NS = SOFTMAX_LOOP_1_C_0;
        end
        else begin
          state_var_NS = CM_LOOP_1_C_0;
        end
      end
      SOFTMAX_LOOP_1_C_0 : begin
        fsm_output = 9'b010101010;
        state_var_NS = SOFTMAX_LOOP_3_C_0;
      end
      SOFTMAX_LOOP_3_C_0 : begin
        fsm_output = 9'b010101011;
        if ( SOFTMAX_LOOP_3_C_0_tr0 ) begin
          state_var_NS = SOFTMAX_LOOP_4_C_0;
        end
        else begin
          state_var_NS = SOFTMAX_LOOP_3_C_0;
        end
      end
      SOFTMAX_LOOP_4_C_0 : begin
        fsm_output = 9'b010101100;
        state_var_NS = SOFTMAX_LOOP_4_C_1;
      end
      SOFTMAX_LOOP_4_C_1 : begin
        fsm_output = 9'b010101101;
        state_var_NS = SOFTMAX_LOOP_4_C_2;
      end
      SOFTMAX_LOOP_4_C_2 : begin
        fsm_output = 9'b010101110;
        if ( SOFTMAX_LOOP_4_C_2_tr0 ) begin
          state_var_NS = SOFTMAX_LOOP_5_C_0;
        end
        else begin
          state_var_NS = SOFTMAX_LOOP_4_C_0;
        end
      end
      SOFTMAX_LOOP_5_C_0 : begin
        fsm_output = 9'b010101111;
        state_var_NS = SOFTMAX_LOOP_5_C_1;
      end
      SOFTMAX_LOOP_5_C_1 : begin
        fsm_output = 9'b010110000;
        state_var_NS = SOFTMAX_LOOP_5_C_2;
      end
      SOFTMAX_LOOP_5_C_2 : begin
        fsm_output = 9'b010110001;
        state_var_NS = SOFTMAX_LOOP_5_C_3;
      end
      SOFTMAX_LOOP_5_C_3 : begin
        fsm_output = 9'b010110010;
        state_var_NS = SOFTMAX_LOOP_5_C_4;
      end
      SOFTMAX_LOOP_5_C_4 : begin
        fsm_output = 9'b010110011;
        state_var_NS = SOFTMAX_LOOP_5_C_5;
      end
      SOFTMAX_LOOP_5_C_5 : begin
        fsm_output = 9'b010110100;
        state_var_NS = SOFTMAX_LOOP_5_C_6;
      end
      SOFTMAX_LOOP_5_C_6 : begin
        fsm_output = 9'b010110101;
        state_var_NS = SOFTMAX_LOOP_5_C_7;
      end
      SOFTMAX_LOOP_5_C_7 : begin
        fsm_output = 9'b010110110;
        state_var_NS = SOFTMAX_LOOP_5_C_8;
      end
      SOFTMAX_LOOP_5_C_8 : begin
        fsm_output = 9'b010110111;
        state_var_NS = SOFTMAX_LOOP_5_C_9;
      end
      SOFTMAX_LOOP_5_C_9 : begin
        fsm_output = 9'b010111000;
        state_var_NS = SOFTMAX_LOOP_5_C_10;
      end
      SOFTMAX_LOOP_5_C_10 : begin
        fsm_output = 9'b010111001;
        state_var_NS = SOFTMAX_LOOP_5_C_11;
      end
      SOFTMAX_LOOP_5_C_11 : begin
        fsm_output = 9'b010111010;
        state_var_NS = SOFTMAX_LOOP_5_C_12;
      end
      SOFTMAX_LOOP_5_C_12 : begin
        fsm_output = 9'b010111011;
        state_var_NS = SOFTMAX_LOOP_5_C_13;
      end
      SOFTMAX_LOOP_5_C_13 : begin
        fsm_output = 9'b010111100;
        state_var_NS = SOFTMAX_LOOP_5_C_14;
      end
      SOFTMAX_LOOP_5_C_14 : begin
        fsm_output = 9'b010111101;
        state_var_NS = SOFTMAX_LOOP_5_C_15;
      end
      SOFTMAX_LOOP_5_C_15 : begin
        fsm_output = 9'b010111110;
        state_var_NS = SOFTMAX_LOOP_5_C_16;
      end
      SOFTMAX_LOOP_5_C_16 : begin
        fsm_output = 9'b010111111;
        state_var_NS = SOFTMAX_LOOP_5_C_17;
      end
      SOFTMAX_LOOP_5_C_17 : begin
        fsm_output = 9'b011000000;
        state_var_NS = SOFTMAX_LOOP_5_C_18;
      end
      SOFTMAX_LOOP_5_C_18 : begin
        fsm_output = 9'b011000001;
        state_var_NS = SOFTMAX_LOOP_5_C_19;
      end
      SOFTMAX_LOOP_5_C_19 : begin
        fsm_output = 9'b011000010;
        if ( SOFTMAX_LOOP_5_C_19_tr0 ) begin
          state_var_NS = SOFTMAX_LOOP_1_C_1;
        end
        else begin
          state_var_NS = SOFTMAX_LOOP_5_C_0;
        end
      end
      SOFTMAX_LOOP_1_C_1 : begin
        fsm_output = 9'b011000011;
        if ( SOFTMAX_LOOP_1_C_1_tr0 ) begin
          state_var_NS = GEMM_3D_FLOAT_LOOP_3_1_C_0;
        end
        else begin
          state_var_NS = SOFTMAX_LOOP_1_C_0;
        end
      end
      GEMM_3D_FLOAT_LOOP_3_1_C_0 : begin
        fsm_output = 9'b011000100;
        state_var_NS = GEMM_3D_FLOAT_LOOP_4_1_C_0;
      end
      GEMM_3D_FLOAT_LOOP_4_1_C_0 : begin
        fsm_output = 9'b011000101;
        state_var_NS = GEMM_3D_FLOAT_LOOP_4_1_C_1;
      end
      GEMM_3D_FLOAT_LOOP_4_1_C_1 : begin
        fsm_output = 9'b011000110;
        state_var_NS = GEMM_3D_FLOAT_LOOP_4_1_C_2;
      end
      GEMM_3D_FLOAT_LOOP_4_1_C_2 : begin
        fsm_output = 9'b011000111;
        state_var_NS = GEMM_3D_FLOAT_LOOP_4_1_C_3;
      end
      GEMM_3D_FLOAT_LOOP_4_1_C_3 : begin
        fsm_output = 9'b011001000;
        if ( GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0 ) begin
          state_var_NS = GEMM_3D_FLOAT_LOOP_3_1_C_1;
        end
        else begin
          state_var_NS = GEMM_3D_FLOAT_LOOP_4_1_C_0;
        end
      end
      GEMM_3D_FLOAT_LOOP_3_1_C_1 : begin
        fsm_output = 9'b011001001;
        if ( GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0 ) begin
          state_var_NS = GEMM_3D_FLOAT_LOOP_1_1_C_0;
        end
        else begin
          state_var_NS = GEMM_3D_FLOAT_LOOP_3_1_C_0;
        end
      end
      GEMM_3D_FLOAT_LOOP_1_1_C_0 : begin
        fsm_output = 9'b011001010;
        if ( GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0 ) begin
          state_var_NS = ATTN_2D_LOOP_3_C_0;
        end
        else begin
          state_var_NS = GEMM_3D_FLOAT_LOOP_3_1_C_0;
        end
      end
      ATTN_2D_LOOP_3_C_0 : begin
        fsm_output = 9'b011001011;
        if ( ATTN_2D_LOOP_3_C_0_tr0 ) begin
          state_var_NS = ATTN_2D_LOOP_2_C_0;
        end
        else begin
          state_var_NS = ATTN_2D_LOOP_3_C_0;
        end
      end
      ATTN_2D_LOOP_2_C_0 : begin
        fsm_output = 9'b011001100;
        if ( ATTN_2D_LOOP_2_C_0_tr0 ) begin
          state_var_NS = RMS_NORM_LOOP_1_2_C_0;
        end
        else begin
          state_var_NS = ATTN_2D_LOOP_3_C_0;
        end
      end
      RMS_NORM_LOOP_1_2_C_0 : begin
        fsm_output = 9'b011001101;
        state_var_NS = RMS_NORM_LOOP_1_2_C_1;
      end
      RMS_NORM_LOOP_1_2_C_1 : begin
        fsm_output = 9'b011001110;
        state_var_NS = RMS_NORM_LOOP_1_2_C_2;
      end
      RMS_NORM_LOOP_1_2_C_2 : begin
        fsm_output = 9'b011001111;
        if ( RMS_NORM_LOOP_1_2_C_2_tr0 ) begin
          state_var_NS = main_C_49;
        end
        else begin
          state_var_NS = RMS_NORM_LOOP_1_2_C_0;
        end
      end
      main_C_49 : begin
        fsm_output = 9'b011010000;
        state_var_NS = compute_sqrt_1_for_C_0;
      end
      compute_sqrt_1_for_C_0 : begin
        fsm_output = 9'b011010001;
        state_var_NS = compute_sqrt_1_for_C_1;
      end
      compute_sqrt_1_for_C_1 : begin
        fsm_output = 9'b011010010;
        state_var_NS = compute_sqrt_1_for_C_2;
      end
      compute_sqrt_1_for_C_2 : begin
        fsm_output = 9'b011010011;
        state_var_NS = compute_sqrt_1_for_C_3;
      end
      compute_sqrt_1_for_C_3 : begin
        fsm_output = 9'b011010100;
        state_var_NS = compute_sqrt_1_for_C_4;
      end
      compute_sqrt_1_for_C_4 : begin
        fsm_output = 9'b011010101;
        state_var_NS = compute_sqrt_1_for_C_5;
      end
      compute_sqrt_1_for_C_5 : begin
        fsm_output = 9'b011010110;
        state_var_NS = compute_sqrt_1_for_C_6;
      end
      compute_sqrt_1_for_C_6 : begin
        fsm_output = 9'b011010111;
        state_var_NS = compute_sqrt_1_for_C_7;
      end
      compute_sqrt_1_for_C_7 : begin
        fsm_output = 9'b011011000;
        state_var_NS = compute_sqrt_1_for_C_8;
      end
      compute_sqrt_1_for_C_8 : begin
        fsm_output = 9'b011011001;
        state_var_NS = compute_sqrt_1_for_C_9;
      end
      compute_sqrt_1_for_C_9 : begin
        fsm_output = 9'b011011010;
        state_var_NS = compute_sqrt_1_for_C_10;
      end
      compute_sqrt_1_for_C_10 : begin
        fsm_output = 9'b011011011;
        state_var_NS = compute_sqrt_1_for_C_11;
      end
      compute_sqrt_1_for_C_11 : begin
        fsm_output = 9'b011011100;
        state_var_NS = compute_sqrt_1_for_C_12;
      end
      compute_sqrt_1_for_C_12 : begin
        fsm_output = 9'b011011101;
        state_var_NS = compute_sqrt_1_for_C_13;
      end
      compute_sqrt_1_for_C_13 : begin
        fsm_output = 9'b011011110;
        state_var_NS = compute_sqrt_1_for_C_14;
      end
      compute_sqrt_1_for_C_14 : begin
        fsm_output = 9'b011011111;
        state_var_NS = compute_sqrt_1_for_C_15;
      end
      compute_sqrt_1_for_C_15 : begin
        fsm_output = 9'b011100000;
        if ( compute_sqrt_1_for_C_15_tr0 ) begin
          state_var_NS = main_C_50;
        end
        else begin
          state_var_NS = compute_sqrt_1_for_C_0;
        end
      end
      main_C_50 : begin
        fsm_output = 9'b011100001;
        state_var_NS = main_C_51;
      end
      main_C_51 : begin
        fsm_output = 9'b011100010;
        state_var_NS = main_C_52;
      end
      main_C_52 : begin
        fsm_output = 9'b011100011;
        state_var_NS = main_C_53;
      end
      main_C_53 : begin
        fsm_output = 9'b011100100;
        state_var_NS = main_C_54;
      end
      main_C_54 : begin
        fsm_output = 9'b011100101;
        state_var_NS = main_C_55;
      end
      main_C_55 : begin
        fsm_output = 9'b011100110;
        state_var_NS = main_C_56;
      end
      main_C_56 : begin
        fsm_output = 9'b011100111;
        state_var_NS = main_C_57;
      end
      main_C_57 : begin
        fsm_output = 9'b011101000;
        state_var_NS = main_C_58;
      end
      main_C_58 : begin
        fsm_output = 9'b011101001;
        state_var_NS = main_C_59;
      end
      main_C_59 : begin
        fsm_output = 9'b011101010;
        state_var_NS = main_C_60;
      end
      main_C_60 : begin
        fsm_output = 9'b011101011;
        state_var_NS = main_C_61;
      end
      main_C_61 : begin
        fsm_output = 9'b011101100;
        state_var_NS = main_C_62;
      end
      main_C_62 : begin
        fsm_output = 9'b011101101;
        state_var_NS = main_C_63;
      end
      main_C_63 : begin
        fsm_output = 9'b011101110;
        state_var_NS = main_C_64;
      end
      main_C_64 : begin
        fsm_output = 9'b011101111;
        state_var_NS = main_C_65;
      end
      main_C_65 : begin
        fsm_output = 9'b011110000;
        state_var_NS = main_C_66;
      end
      main_C_66 : begin
        fsm_output = 9'b011110001;
        state_var_NS = main_C_67;
      end
      main_C_67 : begin
        fsm_output = 9'b011110010;
        state_var_NS = main_C_68;
      end
      main_C_68 : begin
        fsm_output = 9'b011110011;
        state_var_NS = RMS_NORM_LOOP_2_2_C_0;
      end
      RMS_NORM_LOOP_2_2_C_0 : begin
        fsm_output = 9'b011110100;
        state_var_NS = RMS_NORM_LOOP_2_2_C_1;
      end
      RMS_NORM_LOOP_2_2_C_1 : begin
        fsm_output = 9'b011110101;
        state_var_NS = RMS_NORM_LOOP_2_2_C_2;
      end
      RMS_NORM_LOOP_2_2_C_2 : begin
        fsm_output = 9'b011110110;
        state_var_NS = RMS_NORM_LOOP_2_2_C_3;
      end
      RMS_NORM_LOOP_2_2_C_3 : begin
        fsm_output = 9'b011110111;
        state_var_NS = RMS_NORM_LOOP_2_2_C_4;
      end
      RMS_NORM_LOOP_2_2_C_4 : begin
        fsm_output = 9'b011111000;
        if ( RMS_NORM_LOOP_2_2_C_4_tr0 ) begin
          state_var_NS = main_C_69;
        end
        else begin
          state_var_NS = RMS_NORM_LOOP_2_2_C_0;
        end
      end
      main_C_69 : begin
        fsm_output = 9'b011111001;
        state_var_NS = main_C_70;
      end
      main_C_70 : begin
        fsm_output = 9'b011111010;
        state_var_NS = main_C_71;
      end
      main_C_71 : begin
        fsm_output = 9'b011111011;
        state_var_NS = main_C_72;
      end
      main_C_72 : begin
        fsm_output = 9'b011111100;
        state_var_NS = main_C_73;
      end
      main_C_73 : begin
        fsm_output = 9'b011111101;
        state_var_NS = main_C_74;
      end
      main_C_74 : begin
        fsm_output = 9'b011111110;
        state_var_NS = main_C_75;
      end
      main_C_75 : begin
        fsm_output = 9'b011111111;
        state_var_NS = main_C_76;
      end
      main_C_76 : begin
        fsm_output = 9'b100000000;
        state_var_NS = main_C_77;
      end
      main_C_77 : begin
        fsm_output = 9'b100000001;
        state_var_NS = main_C_78;
      end
      main_C_78 : begin
        fsm_output = 9'b100000010;
        state_var_NS = main_C_79;
      end
      main_C_79 : begin
        fsm_output = 9'b100000011;
        state_var_NS = main_C_80;
      end
      main_C_80 : begin
        fsm_output = 9'b100000100;
        state_var_NS = main_C_81;
      end
      main_C_81 : begin
        fsm_output = 9'b100000101;
        state_var_NS = main_C_82;
      end
      main_C_82 : begin
        fsm_output = 9'b100000110;
        state_var_NS = main_C_83;
      end
      main_C_83 : begin
        fsm_output = 9'b100000111;
        state_var_NS = main_C_84;
      end
      main_C_84 : begin
        fsm_output = 9'b100001000;
        state_var_NS = main_C_85;
      end
      main_C_85 : begin
        fsm_output = 9'b100001001;
        state_var_NS = main_C_86;
      end
      main_C_86 : begin
        fsm_output = 9'b100001010;
        state_var_NS = main_C_87;
      end
      main_C_87 : begin
        fsm_output = 9'b100001011;
        state_var_NS = main_C_88;
      end
      main_C_88 : begin
        fsm_output = 9'b100001100;
        state_var_NS = main_C_89;
      end
      main_C_89 : begin
        fsm_output = 9'b100001101;
        state_var_NS = main_C_90;
      end
      main_C_90 : begin
        fsm_output = 9'b100001110;
        state_var_NS = main_C_91;
      end
      main_C_91 : begin
        fsm_output = 9'b100001111;
        state_var_NS = main_C_92;
      end
      main_C_92 : begin
        fsm_output = 9'b100010000;
        state_var_NS = main_C_93;
      end
      main_C_93 : begin
        fsm_output = 9'b100010001;
        state_var_NS = main_C_94;
      end
      main_C_94 : begin
        fsm_output = 9'b100010010;
        state_var_NS = main_C_95;
      end
      main_C_95 : begin
        fsm_output = 9'b100010011;
        state_var_NS = main_C_96;
      end
      main_C_96 : begin
        fsm_output = 9'b100010100;
        state_var_NS = main_C_97;
      end
      main_C_97 : begin
        fsm_output = 9'b100010101;
        state_var_NS = main_C_98;
      end
      main_C_98 : begin
        fsm_output = 9'b100010110;
        state_var_NS = main_C_99;
      end
      main_C_99 : begin
        fsm_output = 9'b100010111;
        state_var_NS = main_C_100;
      end
      main_C_100 : begin
        fsm_output = 9'b100011000;
        state_var_NS = QUANTIZE_ACTIVATION_LOOP_3_1_C_0;
      end
      QUANTIZE_ACTIVATION_LOOP_3_1_C_0 : begin
        fsm_output = 9'b100011001;
        state_var_NS = QUANTIZE_ACTIVATION_LOOP_3_1_C_1;
      end
      QUANTIZE_ACTIVATION_LOOP_3_1_C_1 : begin
        fsm_output = 9'b100011010;
        state_var_NS = QUANTIZE_ACTIVATION_LOOP_3_1_C_2;
      end
      QUANTIZE_ACTIVATION_LOOP_3_1_C_2 : begin
        fsm_output = 9'b100011011;
        if ( QUANTIZE_ACTIVATION_LOOP_3_1_C_2_tr0 ) begin
          state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_0;
        end
        else begin
          state_var_NS = QUANTIZE_ACTIVATION_LOOP_3_1_C_0;
        end
      end
      LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_0 : begin
        fsm_output = 9'b100011100;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0 : begin
        fsm_output = 9'b100011101;
        if ( LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0 ) begin
          state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1;
        end
        else begin
          state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0;
        end
      end
      LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1 : begin
        fsm_output = 9'b100011110;
        if ( LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0 ) begin
          state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_0;
        end
        else begin
          state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_0;
        end
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_0 : begin
        fsm_output = 9'b100011111;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_1;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_1 : begin
        fsm_output = 9'b100100000;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_2;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_2 : begin
        fsm_output = 9'b100100001;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_3;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_3 : begin
        fsm_output = 9'b100100010;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_4;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_4 : begin
        fsm_output = 9'b100100011;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_5;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_5 : begin
        fsm_output = 9'b100100100;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_6;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_6 : begin
        fsm_output = 9'b100100101;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_7;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_7 : begin
        fsm_output = 9'b100100110;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_8;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_8 : begin
        fsm_output = 9'b100100111;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_9;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_9 : begin
        fsm_output = 9'b100101000;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_10;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_10 : begin
        fsm_output = 9'b100101001;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_11;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_11 : begin
        fsm_output = 9'b100101010;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_12;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_12 : begin
        fsm_output = 9'b100101011;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_13;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_13 : begin
        fsm_output = 9'b100101100;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_14;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_14 : begin
        fsm_output = 9'b100101101;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_15;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_15 : begin
        fsm_output = 9'b100101110;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_16;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_16 : begin
        fsm_output = 9'b100101111;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_17;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_17 : begin
        fsm_output = 9'b100110000;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_18;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_18 : begin
        fsm_output = 9'b100110001;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_19;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_19 : begin
        fsm_output = 9'b100110010;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_20;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_20 : begin
        fsm_output = 9'b100110011;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_21;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_21 : begin
        fsm_output = 9'b100110100;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_22;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_22 : begin
        fsm_output = 9'b100110101;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_23;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_23 : begin
        fsm_output = 9'b100110110;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_24;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_24 : begin
        fsm_output = 9'b100110111;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_25;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_25 : begin
        fsm_output = 9'b100111000;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_26;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_26 : begin
        fsm_output = 9'b100111001;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_27;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_27 : begin
        fsm_output = 9'b100111010;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_28;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_28 : begin
        fsm_output = 9'b100111011;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_29;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_29 : begin
        fsm_output = 9'b100111100;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_30;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_30 : begin
        fsm_output = 9'b100111101;
        state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31;
      end
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31 : begin
        fsm_output = 9'b100111110;
        if ( LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31_tr0 ) begin
          state_var_NS = for_1_for_C_0;
        end
        else begin
          state_var_NS = LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_0;
        end
      end
      for_1_for_C_0 : begin
        fsm_output = 9'b100111111;
        state_var_NS = for_1_for_C_1;
      end
      for_1_for_C_1 : begin
        fsm_output = 9'b101000000;
        if ( for_1_for_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = for_1_for_C_0;
        end
      end
      // main_C_0
      default : begin
        fsm_output = 9'b000000000;
        state_var_NS = for_for_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    dut_core_wait_dp
// ------------------------------------------------------------------


module dut_core_wait_dp (
  clk, rst, rms_norm_16_div_cmp_z, core_wen1, rms_norm_16_div_cmp_z_oreg
);
  input clk;
  input rst;
  input [71:0] rms_norm_16_div_cmp_z;
  input core_wen1;
  output [39:0] rms_norm_16_div_cmp_z_oreg;


  // Interconnect Declarations
  reg [39:0] rms_norm_16_div_cmp_z_oreg_pconst_39_0;


  // Interconnect Declarations for Component Instantiations 
  assign rms_norm_16_div_cmp_z_oreg = rms_norm_16_div_cmp_z_oreg_pconst_39_0;
  always @(posedge clk) begin
    if ( rst ) begin
      rms_norm_16_div_cmp_z_oreg_pconst_39_0 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( core_wen1 ) begin
      rms_norm_16_div_cmp_z_oreg_pconst_39_0 <= rms_norm_16_div_cmp_z[39:0];
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dut_core_staller
// ------------------------------------------------------------------


module dut_core_staller (
  en, core_wen1, strm_in_rsci_wen_comp, strm_out_rsci_wen_comp, attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
);
  input en;
  output core_wen1;
  input strm_in_rsci_wen_comp;
  input strm_out_rsci_wen_comp;
  output attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1;



  // Interconnect Declarations for Component Instantiations 
  assign attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 = core_wen1 & en;
  assign core_wen1 = strm_in_rsci_wen_comp & strm_out_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dut_core_strm_out_rsci_strm_out_wait_ctrl
// ------------------------------------------------------------------


module dut_core_strm_out_rsci_strm_out_wait_ctrl (
  strm_out_rsci_iswt0, strm_out_rsci_biwt, strm_out_rsci_irdy
);
  input strm_out_rsci_iswt0;
  output strm_out_rsci_biwt;
  input strm_out_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign strm_out_rsci_biwt = strm_out_rsci_iswt0 & strm_out_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dut_core_strm_in_rsci_strm_in_wait_ctrl
// ------------------------------------------------------------------


module dut_core_strm_in_rsci_strm_in_wait_ctrl (
  strm_in_rsci_iswt0, strm_in_rsci_biwt, strm_in_rsci_ivld
);
  input strm_in_rsci_iswt0;
  output strm_in_rsci_biwt;
  input strm_in_rsci_ivld;



  // Interconnect Declarations for Component Instantiations 
  assign strm_in_rsci_biwt = strm_in_rsci_iswt0 & strm_in_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dut_core_strm_out_rsci
// ------------------------------------------------------------------


module dut_core_strm_out_rsci (
  strm_out_rsc_dat, strm_out_rsc_vld, strm_out_rsc_rdy, strm_out_rsci_oswt, strm_out_rsci_wen_comp,
      strm_out_rsci_idat
);
  output [31:0] strm_out_rsc_dat;
  output strm_out_rsc_vld;
  input strm_out_rsc_rdy;
  input strm_out_rsci_oswt;
  output strm_out_rsci_wen_comp;
  input [31:0] strm_out_rsci_idat;


  // Interconnect Declarations
  wire strm_out_rsci_biwt;
  wire strm_out_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_strm_out_rsci_idat;
  assign nl_strm_out_rsci_idat = {(strm_out_rsci_idat[31:2]) , 2'b00};
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd32)) strm_out_rsci (
      .irdy(strm_out_rsci_irdy),
      .ivld(strm_out_rsci_oswt),
      .idat(nl_strm_out_rsci_idat[31:0]),
      .rdy(strm_out_rsc_rdy),
      .vld(strm_out_rsc_vld),
      .dat(strm_out_rsc_dat)
    );
  dut_core_strm_out_rsci_strm_out_wait_ctrl dut_core_strm_out_rsci_strm_out_wait_ctrl_inst
      (
      .strm_out_rsci_iswt0(strm_out_rsci_oswt),
      .strm_out_rsci_biwt(strm_out_rsci_biwt),
      .strm_out_rsci_irdy(strm_out_rsci_irdy)
    );
  assign strm_out_rsci_wen_comp = (~ strm_out_rsci_oswt) | strm_out_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dut_core_strm_in_rsci
// ------------------------------------------------------------------


module dut_core_strm_in_rsci (
  strm_in_rsc_dat, strm_in_rsc_vld, strm_in_rsc_rdy, strm_in_rsci_oswt, strm_in_rsci_wen_comp,
      strm_in_rsci_idat_mxwt
);
  input [31:0] strm_in_rsc_dat;
  input strm_in_rsc_vld;
  output strm_in_rsc_rdy;
  input strm_in_rsci_oswt;
  output strm_in_rsci_wen_comp;
  output [29:0] strm_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire strm_in_rsci_biwt;
  wire strm_in_rsci_ivld;
  wire [31:0] strm_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd32)) strm_in_rsci (
      .rdy(strm_in_rsc_rdy),
      .vld(strm_in_rsc_vld),
      .dat(strm_in_rsc_dat),
      .irdy(strm_in_rsci_oswt),
      .ivld(strm_in_rsci_ivld),
      .idat(strm_in_rsci_idat)
    );
  dut_core_strm_in_rsci_strm_in_wait_ctrl dut_core_strm_in_rsci_strm_in_wait_ctrl_inst
      (
      .strm_in_rsci_iswt0(strm_in_rsci_oswt),
      .strm_in_rsci_biwt(strm_in_rsci_biwt),
      .strm_in_rsci_ivld(strm_in_rsci_ivld)
    );
  assign strm_in_rsci_idat_mxwt = strm_in_rsci_idat[31:2];
  assign strm_in_rsci_wen_comp = (~ strm_in_rsci_oswt) | strm_in_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dut_core
// ------------------------------------------------------------------


module dut_core (
  clk, en, rst, strm_in_rsc_dat, strm_in_rsc_vld, strm_in_rsc_rdy, strm_out_rsc_dat,
      strm_out_rsc_vld, strm_out_rsc_rdy, attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d,
      attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d, attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d,
      attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d, attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d,
      attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d, attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d,
      attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d, attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d,
      attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d, attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d,
      rms_norm_16_div_cmp_a, rms_norm_16_div_cmp_b, rms_norm_16_div_cmp_z, attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_pff,
      attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_pff, attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_pff,
      attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_pff, attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_pff
);
  input clk;
  input en;
  input rst;
  input [31:0] strm_in_rsc_dat;
  input strm_in_rsc_vld;
  output strm_in_rsc_rdy;
  output [31:0] strm_out_rsc_dat;
  output strm_out_rsc_vld;
  input strm_out_rsc_rdy;
  output attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d;
  output [39:0] attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d;
  output [5:0] attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d;
  output [5:0] attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d;
  output [39:0] attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d;
  input [39:0] attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d;
  output [5:0] attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d;
  output [5:0] attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d;
  input [39:0] attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d;
  output [5:0] attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d;
  output [5:0] attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d;
  output [71:0] rms_norm_16_div_cmp_a;
  output [60:0] rms_norm_16_div_cmp_b;
  input [71:0] rms_norm_16_div_cmp_z;
  output attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_pff;
  output attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_pff;
  output attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_pff;
  output attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_pff;
  output attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_pff;


  // Interconnect Declarations
  wire core_wen1;
  wire strm_in_rsci_wen_comp;
  wire [29:0] strm_in_rsci_idat_mxwt;
  wire strm_out_rsci_wen_comp;
  wire attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1;
  wire [55:0] SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z;
  wire [71:0] LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z;
  wire [39:0] rms_norm_16_div_cmp_z_oreg;
  wire [39:0] operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z;
  reg [23:0] LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_71_48;
  reg [13:0] strm_out_rsci_idat_31_18;
  wire [8:0] fsm_output;
  wire [4:0] RMS_NORM_LOOP_2_2_acc_1_tmp;
  wire [5:0] nl_RMS_NORM_LOOP_2_2_acc_1_tmp;
  wire [2:0] CM_LOOP_3_acc_tmp;
  wire [3:0] nl_CM_LOOP_3_acc_tmp;
  wire [2:0] GEMM_3D_FLOAT_LOOP_3_acc_6_tmp;
  wire [3:0] nl_GEMM_3D_FLOAT_LOOP_3_acc_6_tmp;
  wire CACHE_UPDATE_LOOP_1_and_tmp;
  wire [4:0] LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp;
  wire [5:0] nl_LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp;
  wire for_for_and_tmp;
  wire or_dcpl_4;
  wire and_dcpl;
  wire and_dcpl_1;
  wire or_tmp_11;
  wire or_tmp_48;
  wire or_dcpl_45;
  wire or_dcpl_47;
  wire or_dcpl_54;
  wire or_dcpl_60;
  wire or_dcpl_68;
  wire or_dcpl_79;
  wire or_dcpl_96;
  wire or_tmp_104;
  wire mux_tmp_87;
  wire mux_tmp_91;
  wire nor_tmp_28;
  wire mux_tmp_121;
  wire and_dcpl_26;
  wire and_dcpl_45;
  wire nor_tmp_99;
  wire and_dcpl_57;
  wire and_dcpl_61;
  wire and_dcpl_65;
  wire or_dcpl_332;
  wire or_dcpl_337;
  wire or_dcpl_342;
  wire or_dcpl_351;
  wire or_dcpl_377;
  wire or_tmp_330;
  wire nor_tmp_117;
  wire mux_tmp_363;
  wire not_tmp_253;
  wire or_dcpl_508;
  wire or_dcpl_512;
  wire or_dcpl_584;
  wire or_tmp_464;
  wire or_dcpl_672;
  wire or_tmp_507;
  wire mux_tmp_604;
  wire or_tmp_611;
  wire or_dcpl_770;
  wire or_dcpl_774;
  wire or_dcpl_791;
  wire or_dcpl_794;
  wire and_dcpl_148;
  wire or_tmp_682;
  wire or_dcpl_959;
  wire or_dcpl_961;
  wire and_dcpl_181;
  wire and_dcpl_182;
  wire and_dcpl_185;
  wire and_dcpl_186;
  wire and_dcpl_187;
  wire and_dcpl_189;
  wire and_dcpl_190;
  wire and_dcpl_191;
  wire and_dcpl_192;
  wire and_dcpl_193;
  wire and_dcpl_194;
  wire and_dcpl_197;
  wire and_dcpl_198;
  wire and_dcpl_199;
  wire and_dcpl_200;
  wire and_dcpl_201;
  wire and_dcpl_202;
  wire and_dcpl_203;
  wire and_dcpl_204;
  wire or_dcpl_980;
  wire or_dcpl_983;
  wire or_dcpl_985;
  wire or_dcpl_987;
  wire or_dcpl_988;
  wire or_dcpl_989;
  wire or_dcpl_990;
  wire or_dcpl_991;
  wire or_dcpl_993;
  wire or_dcpl_995;
  wire or_dcpl_996;
  wire or_dcpl_997;
  wire or_dcpl_998;
  wire or_dcpl_999;
  wire or_dcpl_1000;
  wire and_dcpl_205;
  wire and_dcpl_206;
  wire and_dcpl_207;
  wire or_dcpl_1001;
  wire or_dcpl_1002;
  wire or_dcpl_1003;
  wire or_dcpl_1004;
  wire or_dcpl_1005;
  wire or_dcpl_1006;
  wire or_dcpl_1007;
  wire or_dcpl_1008;
  wire or_dcpl_1009;
  wire or_dcpl_1010;
  wire or_dcpl_1011;
  wire or_dcpl_1012;
  wire or_dcpl_1013;
  wire or_dcpl_1014;
  wire or_dcpl_1015;
  wire or_dcpl_1016;
  wire or_dcpl_1017;
  wire or_dcpl_1018;
  wire or_dcpl_1019;
  wire and_dcpl_209;
  wire and_dcpl_211;
  wire and_dcpl_212;
  wire and_dcpl_213;
  wire nor_tmp_261;
  wire and_dcpl_215;
  wire and_dcpl_216;
  wire mux_tmp_787;
  wire mux_tmp_788;
  wire and_dcpl_220;
  wire and_dcpl_221;
  wire and_dcpl_222;
  wire or_dcpl_1020;
  wire or_dcpl_1021;
  wire or_dcpl_1022;
  wire or_dcpl_1023;
  wire or_dcpl_1024;
  wire and_dcpl_226;
  wire or_tmp_704;
  wire or_tmp_708;
  wire and_dcpl_231;
  wire or_dcpl_1025;
  wire and_dcpl_237;
  wire and_dcpl_239;
  wire and_dcpl_240;
  wire or_dcpl_1026;
  wire or_dcpl_1027;
  wire or_dcpl_1028;
  wire or_dcpl_1029;
  wire or_dcpl_1030;
  wire or_dcpl_1031;
  wire or_dcpl_1032;
  wire or_dcpl_1033;
  wire or_dcpl_1034;
  wire or_dcpl_1035;
  wire or_dcpl_1036;
  wire or_dcpl_1037;
  wire or_dcpl_1038;
  wire or_dcpl_1039;
  wire or_dcpl_1040;
  wire or_dcpl_1041;
  wire or_dcpl_1042;
  wire or_dcpl_1043;
  wire or_dcpl_1044;
  wire or_dcpl_1045;
  wire or_dcpl_1046;
  wire and_dcpl_241;
  wire and_dcpl_242;
  wire and_dcpl_243;
  wire and_dcpl_248;
  wire and_dcpl_252;
  wire and_dcpl_255;
  wire and_dcpl_256;
  wire and_dcpl_257;
  wire and_dcpl_258;
  wire and_dcpl_259;
  wire or_tmp_728;
  wire and_dcpl_260;
  wire mux_tmp_824;
  wire or_dcpl_1048;
  wire and_dcpl_261;
  wire and_dcpl_263;
  wire and_dcpl_264;
  wire and_dcpl_265;
  wire or_dcpl_1050;
  wire and_dcpl_268;
  wire and_dcpl_270;
  wire mux_tmp_834;
  wire mux_tmp_836;
  wire and_dcpl_272;
  wire and_dcpl_275;
  wire and_dcpl_276;
  wire nor_tmp_282;
  wire and_dcpl_278;
  wire and_dcpl_279;
  wire or_tmp_742;
  wire mux_tmp_839;
  wire mux_tmp_841;
  wire nor_tmp_285;
  wire and_dcpl_289;
  wire and_dcpl_290;
  wire and_dcpl_291;
  wire and_dcpl_292;
  wire and_dcpl_293;
  wire and_dcpl_294;
  wire and_dcpl_295;
  wire or_tmp_755;
  wire and_dcpl_298;
  wire and_dcpl_302;
  wire or_tmp_757;
  wire or_tmp_762;
  wire mux_tmp_857;
  wire and_dcpl_304;
  wire nor_tmp_289;
  wire and_dcpl_306;
  wire and_dcpl_307;
  wire and_dcpl_308;
  wire nor_tmp_291;
  wire or_tmp_767;
  wire and_dcpl_310;
  wire and_dcpl_312;
  wire and_dcpl_313;
  wire and_dcpl_315;
  wire and_dcpl_316;
  wire and_dcpl_318;
  wire and_dcpl_319;
  wire and_dcpl_321;
  wire and_dcpl_322;
  wire and_dcpl_327;
  wire and_dcpl_328;
  wire and_dcpl_334;
  wire and_dcpl_335;
  wire and_dcpl_336;
  wire and_dcpl_338;
  wire and_dcpl_339;
  wire and_dcpl_341;
  wire and_dcpl_342;
  wire nor_tmp_307;
  wire and_dcpl_344;
  wire and_dcpl_346;
  wire or_tmp_798;
  wire and_dcpl_348;
  wire and_dcpl_349;
  wire and_dcpl_350;
  wire and_dcpl_351;
  wire and_dcpl_352;
  wire and_dcpl_353;
  wire and_dcpl_354;
  wire and_dcpl_355;
  wire and_dcpl_357;
  wire and_dcpl_360;
  wire or_dcpl_1063;
  wire and_dcpl_362;
  wire and_dcpl_363;
  wire and_dcpl_364;
  wire and_dcpl_374;
  wire or_tmp_805;
  wire mux_tmp_906;
  wire or_tmp_808;
  wire mux_tmp_908;
  wire mux_tmp_910;
  wire or_tmp_812;
  wire mux_tmp_915;
  wire or_tmp_813;
  wire mux_tmp_916;
  wire mux_tmp_919;
  wire or_tmp_814;
  wire mux_tmp_922;
  wire mux_tmp_927;
  wire mux_tmp_936;
  wire mux_tmp_937;
  wire and_dcpl_376;
  wire and_dcpl_377;
  wire and_dcpl_381;
  wire and_dcpl_382;
  wire or_tmp_833;
  wire mux_tmp_960;
  wire mux_tmp_967;
  wire mux_tmp_968;
  wire and_dcpl_383;
  wire mux_tmp_975;
  wire and_dcpl_385;
  wire and_dcpl_386;
  wire and_dcpl_388;
  wire or_tmp_861;
  wire and_dcpl_390;
  wire or_tmp_878;
  wire and_dcpl_410;
  wire and_dcpl_413;
  wire nor_tmp_329;
  wire mux_tmp_1027;
  wire and_dcpl_414;
  wire and_dcpl_415;
  wire or_tmp_913;
  wire or_tmp_914;
  wire and_dcpl_417;
  wire and_dcpl_420;
  wire and_dcpl_421;
  wire and_dcpl_422;
  wire or_dcpl_1067;
  wire and_dcpl_425;
  wire or_tmp_922;
  wire or_tmp_923;
  wire mux_tmp_1044;
  wire or_tmp_930;
  wire mux_tmp_1051;
  wire mux_tmp_1052;
  wire or_tmp_931;
  wire or_dcpl_1068;
  wire and_dcpl_432;
  wire and_dcpl_433;
  wire or_dcpl_1070;
  wire or_dcpl_1071;
  wire and_dcpl_438;
  wire and_dcpl_439;
  wire or_tmp_938;
  wire not_tmp_549;
  wire and_dcpl_442;
  wire and_dcpl_448;
  wire and_dcpl_449;
  wire and_dcpl_452;
  wire and_dcpl_453;
  wire or_dcpl_1073;
  wire and_dcpl_458;
  wire or_dcpl_1076;
  wire and_dcpl_461;
  wire and_dcpl_462;
  wire or_dcpl_1077;
  wire or_dcpl_1079;
  wire and_dcpl_467;
  wire and_dcpl_468;
  wire or_dcpl_1081;
  wire and_dcpl_471;
  wire or_dcpl_1083;
  wire and_dcpl_477;
  wire and_dcpl_478;
  wire or_tmp_992;
  wire mux_tmp_1113;
  wire or_tmp_993;
  wire and_dcpl_480;
  wire or_dcpl_1084;
  wire and_dcpl_486;
  wire or_dcpl_1085;
  wire or_dcpl_1086;
  wire or_dcpl_1087;
  wire or_dcpl_1088;
  wire or_dcpl_1089;
  wire mux_tmp_1120;
  wire and_dcpl_511;
  wire and_dcpl_512;
  wire and_dcpl_513;
  wire or_dcpl_1090;
  wire and_dcpl_524;
  wire mux_tmp_1163;
  wire and_dcpl_525;
  wire and_dcpl_528;
  wire or_dcpl_1091;
  wire or_dcpl_1092;
  wire mux_tmp_1178;
  wire mux_tmp_1179;
  wire mux_tmp_1183;
  wire mux_tmp_1185;
  wire mux_tmp_1187;
  wire or_tmp_1035;
  wire and_dcpl_539;
  wire or_tmp_1051;
  wire mux_tmp_1218;
  wire mux_tmp_1219;
  wire mux_tmp_1229;
  wire mux_tmp_1237;
  wire mux_tmp_1238;
  wire or_tmp_1066;
  wire mux_tmp_1240;
  wire mux_tmp_1245;
  wire mux_tmp_1250;
  wire and_dcpl_548;
  wire and_dcpl_549;
  wire and_dcpl_550;
  wire and_dcpl_551;
  wire and_dcpl_552;
  wire and_dcpl_553;
  wire and_dcpl_554;
  wire and_dcpl_557;
  wire mux_tmp_1281;
  wire and_dcpl_564;
  wire and_dcpl_576;
  wire and_dcpl_577;
  wire and_dcpl_581;
  wire or_tmp_1128;
  wire and_dcpl_583;
  wire or_tmp_1132;
  wire or_dcpl_1104;
  wire and_dcpl_585;
  wire and_dcpl_586;
  wire and_dcpl_587;
  wire and_dcpl_588;
  wire and_dcpl_591;
  wire and_dcpl_592;
  wire and_dcpl_595;
  wire and_dcpl_598;
  wire and_dcpl_601;
  wire and_dcpl_604;
  wire and_dcpl_607;
  wire and_dcpl_610;
  wire and_dcpl_613;
  wire and_dcpl_616;
  wire and_dcpl_618;
  wire and_dcpl_619;
  wire or_tmp_1203;
  wire and_dcpl_620;
  wire mux_tmp_1421;
  wire or_tmp_1218;
  wire not_tmp_650;
  wire and_dcpl_622;
  wire and_dcpl_625;
  wire or_tmp_1221;
  wire mux_tmp_1426;
  wire and_dcpl_626;
  wire and_dcpl_628;
  wire and_dcpl_629;
  wire mux_tmp_1440;
  wire and_dcpl_635;
  wire and_tmp_42;
  wire mux_tmp_1451;
  wire and_dcpl_641;
  wire and_dcpl_642;
  wire or_dcpl_1108;
  wire mux_tmp_1489;
  wire or_dcpl_1109;
  wire or_dcpl_1114;
  wire and_dcpl_650;
  wire and_dcpl_651;
  wire or_dcpl_1116;
  wire and_dcpl_656;
  wire or_dcpl_1118;
  wire or_dcpl_1119;
  wire or_dcpl_1120;
  wire or_dcpl_1121;
  wire or_dcpl_1122;
  wire or_dcpl_1123;
  wire or_dcpl_1125;
  wire or_dcpl_1126;
  wire or_dcpl_1127;
  wire or_dcpl_1128;
  wire or_dcpl_1130;
  wire or_dcpl_1131;
  wire or_dcpl_1132;
  wire or_dcpl_1133;
  wire or_tmp_1291;
  wire or_tmp_1296;
  wire and_dcpl_718;
  wire or_tmp_1316;
  wire mux_tmp_1519;
  wire or_tmp_1320;
  wire and_dcpl_721;
  wire not_tmp_699;
  wire and_dcpl_725;
  wire and_dcpl_726;
  wire or_dcpl_1134;
  wire or_dcpl_1137;
  wire or_dcpl_1138;
  wire or_dcpl_1140;
  wire or_dcpl_1141;
  wire and_dcpl_727;
  wire and_dcpl_728;
  wire and_dcpl_729;
  wire and_dcpl_730;
  wire and_dcpl_731;
  wire and_dcpl_732;
  wire mux_tmp_1548;
  wire mux_tmp_1549;
  wire nand_tmp_66;
  wire and_dcpl_735;
  wire and_dcpl_736;
  wire and_dcpl_739;
  wire and_dcpl_740;
  wire and_dcpl_743;
  wire and_dcpl_745;
  wire and_dcpl_747;
  wire and_dcpl_748;
  wire mux_tmp_1562;
  wire and_dcpl_751;
  wire and_dcpl_753;
  wire and_dcpl_754;
  wire and_dcpl_758;
  wire and_dcpl_760;
  wire and_dcpl_764;
  wire and_dcpl_768;
  wire and_dcpl_772;
  wire and_dcpl_776;
  wire and_dcpl_780;
  wire and_dcpl_784;
  wire and_dcpl_788;
  wire and_dcpl_792;
  wire and_dcpl_796;
  wire and_dcpl_800;
  wire and_dcpl_804;
  wire and_dcpl_810;
  wire and_dcpl_812;
  wire and_dcpl_813;
  wire and_dcpl_814;
  wire mux_tmp_1578;
  wire and_dcpl_817;
  wire and_dcpl_818;
  wire and_dcpl_819;
  wire and_dcpl_820;
  wire and_dcpl_821;
  wire or_tmp_1354;
  wire and_dcpl_825;
  wire and_dcpl_826;
  wire and_dcpl_827;
  wire and_dcpl_830;
  wire and_dcpl_831;
  wire and_dcpl_832;
  wire and_dcpl_835;
  wire and_dcpl_836;
  wire and_dcpl_837;
  wire and_dcpl_840;
  wire and_dcpl_841;
  wire and_dcpl_842;
  wire and_dcpl_843;
  wire and_dcpl_847;
  wire and_dcpl_850;
  wire and_dcpl_851;
  wire and_dcpl_854;
  wire and_dcpl_855;
  wire and_dcpl_856;
  wire and_dcpl_859;
  wire and_dcpl_860;
  wire and_dcpl_863;
  wire and_dcpl_864;
  wire and_dcpl_867;
  wire and_dcpl_868;
  wire and_dcpl_871;
  wire and_dcpl_872;
  wire and_dcpl_875;
  wire and_dcpl_876;
  wire and_dcpl_879;
  wire and_dcpl_880;
  wire and_dcpl_885;
  wire or_tmp_1392;
  wire and_dcpl_888;
  wire and_dcpl_959;
  wire mux_tmp_1943;
  wire mux_tmp_1945;
  wire and_dcpl_983;
  wire and_dcpl_987;
  wire and_dcpl_989;
  wire and_dcpl_999;
  wire and_dcpl_1000;
  wire mux_tmp_1990;
  wire mux_tmp_1993;
  wire and_dcpl_1003;
  wire or_dcpl_1145;
  wire mux_tmp_2013;
  wire mux_tmp_2015;
  wire or_dcpl_1146;
  wire mux_tmp_2034;
  wire and_dcpl_1011;
  wire and_dcpl_1033;
  wire and_dcpl_1034;
  wire mux_tmp_2067;
  wire and_dcpl_1055;
  wire and_dcpl_1061;
  wire or_tmp_1632;
  wire not_tmp_874;
  wire or_tmp_1643;
  wire or_dcpl_1152;
  wire or_dcpl_1155;
  wire or_dcpl_1156;
  wire or_dcpl_1158;
  wire or_dcpl_1159;
  wire or_dcpl_1160;
  wire or_dcpl_1161;
  wire or_dcpl_1162;
  wire or_dcpl_1163;
  wire or_dcpl_1164;
  wire or_dcpl_1165;
  wire or_dcpl_1166;
  wire or_dcpl_1167;
  wire or_dcpl_1168;
  wire or_dcpl_1169;
  wire or_dcpl_1170;
  wire and_dcpl_1073;
  wire and_dcpl_1082;
  wire and_dcpl_1084;
  wire and_dcpl_1088;
  wire and_dcpl_1091;
  wire and_dcpl_1094;
  wire and_dcpl_1097;
  wire and_dcpl_1100;
  wire and_dcpl_1103;
  wire and_dcpl_1106;
  wire and_dcpl_1109;
  wire and_dcpl_1112;
  wire and_dcpl_1115;
  wire and_dcpl_1118;
  wire and_dcpl_1121;
  wire and_dcpl_1124;
  wire and_dcpl_1127;
  wire and_dcpl_1130;
  wire and_dcpl_1141;
  wire and_dcpl_1145;
  wire and_dcpl_1151;
  wire and_dcpl_1152;
  wire or_tmp_1664;
  wire mux_tmp_2116;
  wire nand_tmp_99;
  wire mux_tmp_2119;
  wire or_tmp_1671;
  wire mux_tmp_2121;
  wire and_dcpl_1154;
  wire and_dcpl_1162;
  wire or_tmp_1690;
  wire mux_tmp_2153;
  wire or_dcpl_1178;
  wire mux_tmp_2176;
  wire or_dcpl_1180;
  wire or_dcpl_1181;
  wire or_dcpl_1183;
  wire or_dcpl_1184;
  wire or_dcpl_1186;
  wire or_dcpl_1187;
  wire or_dcpl_1188;
  wire or_dcpl_1189;
  wire and_dcpl_1193;
  wire and_dcpl_1194;
  wire and_dcpl_1195;
  wire or_dcpl_1195;
  wire or_dcpl_1196;
  wire or_dcpl_1198;
  wire or_dcpl_1199;
  wire or_dcpl_1201;
  wire or_dcpl_1203;
  wire or_dcpl_1209;
  wire and_dcpl_1199;
  wire nand_tmp_104;
  wire mux_tmp_2252;
  wire and_dcpl_1225;
  wire and_dcpl_1227;
  wire and_dcpl_1232;
  wire QUANTIZE_ACTIVATION_LOOP_3_nand_seb;
  wire QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse;
  wire RESHAPE_2D_TO_3D_LOOP_2_2_and_cse;
  reg [4:0] RMS_NORM_LOOP_2_2_i_4_0_sva_1;
  reg RMS_NORM_LOOP_2_2_and_30_m1c;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1;
  wire RMS_NORM_LOOP_2_2_and_30_m1c_1;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_2_mx0;
  wire [35:0] operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1;
  wire [36:0] nl_operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1;
  wire GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_1_sva_1;
  wire GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_2_sva_1;
  wire GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_3_sva_1;
  wire GEMM_3D_FLOAT_LOOP_3_and_stg_2_0_sva_1;
  wire GEMM_3D_FLOAT_LOOP_3_and_stg_2_1_sva_1;
  wire GEMM_3D_FLOAT_LOOP_3_and_stg_2_2_sva_1;
  wire GEMM_3D_FLOAT_LOOP_3_and_stg_2_3_sva_1;
  wire GEMM_3D_FLOAT_LOOP_3_and_stg_1_0_sva_1;
  wire GEMM_3D_FLOAT_LOOP_3_and_stg_1_1_sva_1;
  wire GEMM_3D_FLOAT_LOOP_3_and_stg_1_2_sva_1;
  wire GEMM_3D_FLOAT_LOOP_3_and_stg_1_3_sva_1;
  reg RMS_NORM_LOOP_2_and_30_m1c;
  wire RMS_NORM_LOOP_2_and_30_m1c_1;
  reg [4:0] LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1;
  reg GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva;
  reg GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva;
  reg GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva;
  reg GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva;
  reg GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva;
  reg GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva;
  reg GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva;
  reg GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva;
  reg GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva;
  reg GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva;
  reg GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva;
  reg GEMM_3D_FLOAT_LOOP_3_and_tmp_sva;
  reg [39:0] RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva;
  reg [39:0] input_0_0_sva_2;
  reg GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva;
  reg [2:0] TRANSPOSE_LAST_TWO_DIMS_LOOP_3_k_2_0_sva_1;
  reg GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva;
  reg [39:0] RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva;
  wire [1:0] LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_conc_1_1_1_0_svs_1;
  wire RMS_NORM_LOOP_2_2_unequal_tmp_mx0w0;
  wire GEMM_3D_FLOAT_LOOP_4_l_and_ssc;
  reg reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd;
  reg reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  wire and_336_ssc;
  wire mux_856_ssc;
  reg [20:0] LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_59_39;
  reg [38:0] LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_38_0;
  wire mux_851_ssc;
  wire and_321_ssc;
  reg operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_39;
  reg [3:0] operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_38_35;
  wire mux_2100_ssc;
  reg LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1;
  reg LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0;
  wire attention_abs_qelse_and_ssc;
  wire attention_abs_4_qelse_and_ssc;
  wire for_1_for_and_cse;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_and_cse;
  wire input_and_cse;
  wire and_1555_cse;
  wire or_1769_cse;
  wire or_1732_cse;
  wire or_1770_cse;
  reg reg_strm_out_rsci_iswt0_cse;
  reg reg_strm_in_rsci_iswt0_cse;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_and_3_cse;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_and_6_cse;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_and_7_cse;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_and_8_cse;
  wire and_1474_cse;
  wire and_1559_cse;
  wire mux_806_cse;
  wire or_2249_cse;
  wire and_1773_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_cse;
  wire or_2456_cse;
  wire and_1651_cse;
  wire or_1907_cse;
  wire nand_365_cse;
  wire or_2480_cse;
  wire or_2486_cse;
  wire or_2742_cse;
  wire or_2736_cse;
  wire or_1880_cse;
  wire mux_792_cse;
  wire or_1983_cse;
  wire or_2457_cse;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_and_28_cse;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_and_cse;
  wire GEMM_3D_FLOAT_LOOP_3_1_and_44_cse;
  wire [39:0] attention_2_1_16_16_4_4_q_embed_mux_14_cse;
  wire [39:0] attention_2_1_16_16_4_4_q_embed_mux_13_cse;
  wire attention_2_1_16_16_4_4_q_embed_and_cse;
  wire [39:0] attention_2_1_16_16_4_4_q_embed_mux_11_cse;
  wire [39:0] attention_2_1_16_16_4_4_q_embed_mux_9_cse;
  wire [39:0] attention_2_1_16_16_4_4_q_embed_mux_7_cse;
  wire nor_1239_cse;
  wire attention_2_1_16_16_4_4_attn_weights_and_cse;
  wire GEMM_3D_FLOAT_LOOP_3_and_36_cse;
  wire attention_2_1_16_16_4_4_attn_weights_and_12_cse;
  wire attention_2_1_16_16_4_4_attn_weights_and_24_cse;
  wire GEMM_3D_FLOAT_LOOP_3_1_and_46_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_8_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_16_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_24_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_32_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_40_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_48_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_56_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_64_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_72_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_80_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_88_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_96_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_104_cse;
  wire attention_2_1_16_16_4_4_quantized_final_output_and_112_cse;
  wire and_1455_cse;
  wire nor_176_cse;
  wire or_76_cse;
  wire or_130_cse;
  wire and_28_cse;
  wire nor_1229_cse;
  wire and_1771_cse;
  wire and_1762_cse;
  wire or_3185_cse;
  wire nor_366_cse;
  wire nand_197_cse;
  wire or_2699_cse;
  wire or_1848_cse;
  wire or_133_cse;
  wire nor_777_cse;
  wire nor_973_cse;
  wire and_37_cse;
  wire or_361_cse;
  wire or_362_cse;
  wire and_1638_cse;
  wire or_1985_cse;
  wire or_1984_cse;
  wire nor_749_cse;
  wire or_2455_cse;
  wire or_1197_cse;
  wire or_822_cse;
  wire or_2460_cse;
  wire or_1879_cse;
  wire nor_1026_cse;
  wire or_270_cse;
  wire or_1767_cse;
  wire or_1772_cse;
  wire nor_717_cse;
  wire and_1572_cse;
  wire or_1908_cse;
  wire or_255_cse;
  wire or_1851_cse;
  wire or_1835_cse;
  wire or_1867_cse;
  wire or_1420_cse;
  wire mux_623_cse;
  wire mux_528_cse;
  wire and_1570_cse;
  wire or_750_cse;
  wire or_619_cse;
  wire or_790_cse;
  wire nand_143_cse;
  wire or_262_cse;
  wire or_1435_cse;
  wire or_806_cse;
  wire or_1431_cse;
  wire or_753_cse;
  wire nor_992_cse;
  wire or_2792_cse;
  wire or_1795_cse;
  wire nand_253_cse;
  wire or_349_cse;
  wire or_241_cse;
  wire or_2451_cse;
  wire nor_646_cse;
  wire nand_129_cse;
  wire or_3167_cse;
  wire nor_354_cse;
  wire nor_355_cse;
  wire or_2395_cse;
  wire nand_163_cse;
  wire nand_240_cse;
  wire nor_964_cse;
  wire nand_263_cse;
  wire or_2834_cse;
  wire or_2797_cse;
  wire nand_381_cse;
  wire or_2029_cse;
  wire nor_1106_cse;
  wire nor_593_cse;
  wire or_2500_cse;
  wire or_2154_cse;
  wire or_2739_cse;
  wire or_3039_cse;
  wire and_1782_cse;
  wire or_3163_cse;
  wire nor_305_cse;
  wire or_2671_cse;
  wire and_1790_cse;
  wire mux_816_ssc;
  reg reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd;
  reg reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd_1;
  wire RMS_NORM_LOOP_2_2_i_and_ssc;
  reg [2:0] reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd;
  reg reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1;
  reg [23:0] reg_rms_norm_16_div_cmp_a_ftd;
  wire and_937_ssc;
  wire nor_1324_seb;
  wire CACHE_UPDATE_LOOP_3_k_and_ssc;
  reg reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  reg [1:0] operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_17_16;
  reg reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1;
  reg reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0;
  wire for_for_and_13_ssc;
  wire QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_or_cse;
  wire mux_1639_cse;
  wire mux_1551_cse;
  wire or_2481_cse;
  wire mux_1812_cse;
  wire mux_1809_cse;
  wire mux_2025_cse;
  wire mux_2157_cse;
  wire mux_958_cse;
  wire and_1637_cse;
  wire mux_2024_cse;
  wire or_2717_cse;
  wire mux_502_cse;
  wire mux_304_cse;
  wire mux_1522_cse;
  wire or_3137_cse;
  wire mux_624_cse;
  wire nor_998_cse;
  wire nand_50_cse;
  wire mux_1074_cse;
  wire mux_1089_cse;
  wire mux_1087_cse;
  wire mux_1084_cse;
  wire mux_1309_cse;
  wire mux_2092_cse;
  wire and_1811_cse;
  wire and_1781_cse;
  wire mux_2139_cse;
  wire or_2858_cse;
  wire or_2856_cse;
  wire attention_2_1_16_16_4_4_attn_output_and_4_cse;
  wire attention_2_1_16_16_4_4_attn_weights_and_36_cse;
  wire attention_2_1_16_16_4_4_q_embed_and_5_cse;
  wire mux_1559_cse;
  wire mux_1557_cse;
  wire mux_1555_cse;
  wire mux_1553_cse;
  wire mux_1645_cse;
  wire mux_1546_cse;
  wire mux_2032_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_32_cse;
  wire attention_2_1_16_16_4_4_attn_weights_and_48_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_63_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_65_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_67_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_69_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_71_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_73_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_75_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_77_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_79_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_81_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_83_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_85_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_87_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_89_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_91_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_93_cse;
  wire output_and_16_cse;
  wire mux_1122_cse;
  wire mux_1125_cse;
  wire RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c4;
  wire and_1191_rgt;
  wire and_622_rgt;
  wire operator_40_24_true_AC_TRN_AC_WRAP_1_and_ssc;
  reg operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_15;
  wire mux_1132_cse;
  wire [19:0] CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_sdt;
  wire and_362_ssc;
  reg [2:0] TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_16_psp_1;
  wire [3:0] nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_16_psp_1;
  wire [2:0] GEMM_3D_FLOAT_LOOP_4_acc_sdt_1;
  wire [3:0] nl_GEMM_3D_FLOAT_LOOP_4_acc_sdt_1;
  wire [2:0] GEMM_3D_FLOAT_LOOP_4_acc_13_sdt_1;
  wire [3:0] nl_GEMM_3D_FLOAT_LOOP_4_acc_13_sdt_1;
  wire [2:0] GEMM_3D_FLOAT_LOOP_4_1_acc_12_sdt_1;
  wire [3:0] nl_GEMM_3D_FLOAT_LOOP_4_1_acc_12_sdt_1;
  wire [2:0] CACHE_UPDATE_LOOP_3_acc_sdt_1;
  wire [3:0] nl_CACHE_UPDATE_LOOP_3_acc_sdt_1;
  wire [2:0] TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_sdt_1;
  wire [3:0] nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_sdt_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_0_0_0_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_2_0_3_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_3_0_0_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_3_0_1_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_3_0_2_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_15_0;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0;
  wire and_dcpl_1233;
  wire [35:0] attention_abs_qr_35_0_lpi_1_dfm_mx0w0;
  wire [36:0] nl_attention_abs_qr_35_0_lpi_1_dfm_mx0w0;
  wire GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva_mx0w0;
  wire GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva_mx0w0;
  wire GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva_mx0w0;
  wire attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c10;
  reg [39:0] input_0_4_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3;
  wire attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c0;
  wire attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c1;
  wire attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c10;
  reg [39:0] input_0_11_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3;
  wire attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c0;
  wire attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c1;
  wire attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c10;
  reg [39:0] input_0_3_sva_1;
  reg [5:0] for_for_strm_in_tmp_sva_31_26;
  reg [23:0] for_for_strm_in_tmp_sva_25_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3;
  wire attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c0;
  wire attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c1;
  wire attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c12;
  wire or_3212_tmp;
  wire or_3213_tmp;
  wire or_3214_tmp;
  wire nand_303_tmp;
  wire nand_304_tmp;
  wire nand_305_tmp;
  wire and_343_itm;
  wire [39:0] GEMM_3D_FLOAT_LOOP_4_1_mux1h_5_itm;
  wire and_404_itm;
  wire and_416_itm;
  wire and_428_itm;
  wire [7:0] LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_itm;
  wire [7:0] LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_itm;
  wire [14:0] APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_itm;
  wire and_615_itm;
  wire and_633_itm;
  wire and_654_itm;
  wire and_648_itm;
  wire and_642_itm;
  wire and_636_itm;
  wire and_629_itm;
  wire and_639_itm;
  wire and_645_itm;
  wire and_651_itm;
  wire and_657_itm;
  wire nor_1144_itm;
  wire [12:0] APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm;
  wire and_1060_itm;
  wire [7:0] LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm;
  wire [7:0] LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm;
  wire mux_2256_itm;
  wire mux_1147_itm;
  wire mux_1177_itm;
  wire mux_1197_itm;
  wire [18:0] CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_itm;
  wire and_dcpl_1248;
  wire [15:0] z_out;
  wire and_dcpl_1261;
  wire [15:0] z_out_1;
  wire and_dcpl_1273;
  wire [39:0] z_out_2;
  wire and_dcpl_1294;
  wire [2:0] z_out_3;
  wire [3:0] nl_z_out_3;
  wire [2:0] z_out_4;
  wire [3:0] nl_z_out_4;
  wire [2:0] z_out_5;
  wire [3:0] nl_z_out_5;
  wire and_dcpl_1363;
  wire and_dcpl_1371;
  wire and_dcpl_1379;
  wire and_dcpl_1385;
  wire [59:0] z_out_9;
  wire signed [60:0] nl_z_out_9;
  wire and_dcpl_1391;
  wire and_dcpl_1392;
  wire and_dcpl_1393;
  wire and_dcpl_1396;
  wire and_dcpl_1398;
  wire and_dcpl_1401;
  wire and_dcpl_1403;
  wire and_dcpl_1406;
  wire and_dcpl_1407;
  wire and_dcpl_1410;
  wire and_dcpl_1415;
  wire and_dcpl_1420;
  wire and_dcpl_1425;
  wire and_dcpl_1427;
  wire and_dcpl_1429;
  wire and_dcpl_1431;
  wire and_dcpl_1436;
  wire [63:0] z_out_10;
  wire signed [79:0] nl_z_out_10;
  wire and_dcpl_1447;
  wire [2:0] z_out_11;
  wire [3:0] nl_z_out_11;
  wire [4:0] z_out_12;
  wire [5:0] nl_z_out_12;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2;
  reg [39:0] input_0_7_sva_1;
  reg [39:0] input_0_8_sva_1;
  reg [39:0] input_0_6_sva_1;
  reg [39:0] input_0_9_sva_1;
  reg [39:0] input_0_5_sva_1;
  reg [39:0] input_0_10_sva_1;
  reg [39:0] input_0_12_sva_1;
  reg [39:0] input_0_1_sva_1;
  reg [39:0] input_0_14_sva_1;
  reg [39:0] input_0_7_sva_2;
  reg [39:0] input_0_8_sva_2;
  reg [39:0] input_0_6_sva_2;
  reg [39:0] input_0_9_sva_2;
  reg [39:0] input_0_5_sva_2;
  reg [39:0] input_0_10_sva_2;
  reg [39:0] input_0_4_sva_2;
  reg [39:0] input_0_11_sva_2;
  reg [39:0] input_0_3_sva_2;
  reg [39:0] input_0_12_sva_2;
  reg [39:0] input_0_1_sva_2;
  reg [39:0] input_0_14_sva_2;
  reg [39:0] input_0_15_sva_1;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm;
  reg [39:0] apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_2_0_3_lpi_3;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_3_0_0_lpi_3;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_3_0_1_lpi_3;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_3_0_2_lpi_3;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_3_0_3_lpi_3;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_2_0_1_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_1_0_1_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_2_0_3_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_3_0_0_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_0_0_2_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_3_0_1_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_3_0_2_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_0_0_0_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_q_embed_3_0_3_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_4;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_5;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_4;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_4;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_5;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_4;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_4;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_5;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_4;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_4;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_5;
  reg [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_4;
  reg [39:0] softmax_1_4_3_sum_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_3_0_0_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_3_0_1_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_3_0_2_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_3_0_3_sva_2;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1;
  reg [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1;
  reg [39:0] QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva;
  reg RMS_NORM_LOOP_2_and_29_ssc;
  reg RMS_NORM_LOOP_2_and_34_ssc;
  reg RMS_NORM_LOOP_2_2_and_29_ssc;
  reg RMS_NORM_LOOP_2_2_and_34_ssc;
  reg [59:0] LINEAR_FORWARD_NO_MUL_LOOP_2_2_mul_mut;
  reg [59:0] LINEAR_FORWARD_NO_MUL_LOOP_2_3_mul_mut;
  reg [60:0] LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut;
  reg RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_mux1h_itm;
  reg [59:0] LINEAR_FORWARD_NO_MUL_LOOP_2_mul_itm;
  reg [55:0] APPLY_ROTARY_POS_EMB_LOOP_6_mul_itm;
  reg [55:0] APPLY_ROTARY_POS_EMB_LOOP_6_mul_1_itm;
  reg [55:0] APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm;
  reg [55:0] APPLY_ROTARY_POS_EMB_LOOP_6_mul_3_itm;
  wire signed [56:0] nl_APPLY_ROTARY_POS_EMB_LOOP_6_mul_3_itm;
  reg [39:0] GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm;
  reg RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_mux1h_itm;
  reg [38:0] QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_38_0;
  reg [38:0] QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_38_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_7_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_8_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_6_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_9_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_5_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_10_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_4_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_11_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_3_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_12_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_2_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_13_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_1_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_14_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_0_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_re_0_15_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_7_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_8_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_6_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_9_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_5_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_10_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_4_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_11_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_3_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_12_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_2_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_13_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_1_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_14_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_0_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_15_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_7_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_8_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_6_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_9_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_5_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_10_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_4_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_11_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_3_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_12_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_2_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_13_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_1_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_14_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_0_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_15_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_re_0_7_sva_2_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_39_16;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_15_0;
  reg [23:0] attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_39_16;
  reg [15:0] attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_39_16;
  reg [15:0] attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_39_16;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0;
  reg [23:0] attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16;
  reg [15:0] attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16;
  reg [15:0] apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_39_16;
  reg [15:0] apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16;
  reg [23:0] apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16;
  reg [23:0] output_0_7_lpi_3_39_16;
  reg [15:0] output_0_7_lpi_3_15_0;
  reg [23:0] output_0_8_lpi_3_39_16;
  reg [15:0] output_0_8_lpi_3_15_0;
  reg [23:0] output_0_6_lpi_3_39_16;
  reg [15:0] output_0_6_lpi_3_15_0;
  reg [23:0] output_0_9_lpi_3_39_16;
  reg [15:0] output_0_9_lpi_3_15_0;
  reg [23:0] output_0_5_lpi_3_39_16;
  reg [15:0] output_0_5_lpi_3_15_0;
  reg [23:0] output_0_10_lpi_3_39_16;
  reg [15:0] output_0_10_lpi_3_15_0;
  reg [23:0] output_0_4_lpi_3_39_16;
  reg [15:0] output_0_4_lpi_3_15_0;
  reg [23:0] output_0_11_lpi_3_39_16;
  reg [15:0] output_0_11_lpi_3_15_0;
  reg [23:0] output_0_3_lpi_3_39_16;
  reg [15:0] output_0_3_lpi_3_15_0;
  reg [23:0] output_0_12_lpi_3_39_16;
  reg [15:0] output_0_12_lpi_3_15_0;
  reg [23:0] output_0_2_lpi_3_39_16;
  reg [15:0] output_0_2_lpi_3_15_0;
  reg [23:0] output_0_13_lpi_3_39_16;
  reg [15:0] output_0_13_lpi_3_15_0;
  reg [23:0] output_0_1_lpi_3_39_16;
  reg [23:0] output_0_14_lpi_3_39_16;
  reg [15:0] output_0_14_lpi_3_15_0;
  reg [23:0] output_0_0_lpi_3_39_16;
  reg [15:0] output_0_0_lpi_3_15_0;
  reg [23:0] output_0_15_lpi_3_39_16;
  reg [15:0] output_0_15_lpi_3_15_0;
  reg [23:0] output_0_7_lpi_4_39_16;
  reg [23:0] output_0_8_lpi_4_39_16;
  reg [23:0] output_0_6_lpi_4_39_16;
  reg [23:0] output_0_9_lpi_4_39_16;
  reg [23:0] output_0_5_lpi_4_39_16;
  reg [23:0] output_0_10_lpi_4_39_16;
  reg [23:0] output_0_4_lpi_4_39_16;
  reg [23:0] output_0_11_lpi_4_39_16;
  reg [23:0] output_0_3_lpi_4_39_16;
  reg [23:0] output_0_12_lpi_4_39_16;
  reg [23:0] output_0_2_lpi_4_39_16;
  reg [23:0] output_0_13_lpi_4_39_16;
  reg [23:0] output_0_1_lpi_4_39_16;
  reg [23:0] output_0_14_lpi_4_39_16;
  reg [23:0] output_0_0_lpi_4_39_16;
  reg [23:0] output_0_15_lpi_4_39_16;
  reg [23:0] output_0_7_sva_1_39_16;
  reg [23:0] output_0_8_sva_1_39_16;
  reg [23:0] output_0_6_sva_1_39_16;
  reg [23:0] output_0_9_sva_1_39_16;
  reg [23:0] output_0_5_sva_1_39_16;
  reg [23:0] output_0_10_sva_1_39_16;
  reg [23:0] output_0_4_sva_1_39_16;
  reg [23:0] output_0_11_sva_1_39_16;
  reg [23:0] output_0_3_sva_1_39_16;
  reg [23:0] output_0_12_sva_1_39_16;
  reg [23:0] output_0_2_sva_1_39_16;
  reg [23:0] output_0_13_sva_1_39_16;
  reg [23:0] output_0_1_sva_1_39_16;
  reg [23:0] output_0_14_sva_1_39_16;
  reg [23:0] output_0_0_sva_1_39_16;
  reg [23:0] output_0_15_sva_1_39_16;
  reg [15:0] output_0_7_sva_2_15_0;
  reg [15:0] output_0_8_sva_2_15_0;
  reg [15:0] output_0_6_sva_2_15_0;
  reg [15:0] output_0_9_sva_2_15_0;
  reg [15:0] output_0_5_sva_2_15_0;
  reg [15:0] output_0_10_sva_2_15_0;
  reg [15:0] output_0_4_sva_2_15_0;
  reg [15:0] output_0_11_sva_2_15_0;
  reg [15:0] output_0_3_sva_2_15_0;
  reg [15:0] output_0_12_sva_2_15_0;
  reg [15:0] output_0_2_sva_2_15_0;
  reg [15:0] output_0_13_sva_2_15_0;
  reg [15:0] output_0_14_sva_2_15_0;
  reg [15:0] output_0_0_sva_2_15_0;
  reg [15:0] output_0_15_sva_2_15_0;
  reg [23:0] LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48;
  reg [23:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16;
  reg [23:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_39_16;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_7;
  reg attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2_mx1;
  wire [39:0] attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1_mx0w1;
  wire [39:0] attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0_mx0w1;
  wire [39:0] apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2_mx0w1;
  wire [39:0] apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2_mx0w1;
  wire [39:0] apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2_mx0w1;
  wire [39:0] apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2_mx0w1;
  wire [39:0] apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w0;
  wire [39:0] apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w3;
  wire [39:0] apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2_mx0w1;
  wire [23:0] apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16_mx0w1;
  wire [23:0] apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16_mx0w1;
  wire [23:0] apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16_mx0w1;
  wire [23:0] apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16_mx0w1;
  wire [23:0] apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16_mx0w1;
  wire [15:0] attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0_mx0w1;
  wire [15:0] drf_output_sdt_2_sva_15_0_mx0w0;
  wire [15:0] drf_output_sdt_3_sva_15_0_mx0w3;
  wire [39:0] SOFTMAX_LOOP_5_mux_12_psp_mx0w0;
  wire [23:0] LINEAR_FORWARD_NO_MUL_LOOP_2_2_conc_1_mut_71_48_mx0w0;
  wire [23:0] LINEAR_FORWARD_NO_MUL_LOOP_2_3_conc_1_mut_71_48_mx0w3;
  wire [60:0] LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2;
  wire signed [61:0] nl_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2;
  wire rms_norm_16_div_cmp_a_mx0c0;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c0;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c9;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx2;
  wire [39:0] attention_abs_1_qr_sva_1;
  wire [40:0] nl_attention_abs_1_qr_sva_1;
  wire [39:0] softmax_1_4_3_sum_sva_2;
  wire [40:0] nl_softmax_1_4_3_sum_sva_2;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c0;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c2;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c3;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c5;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c7;
  wire for_for_strm_in_tmp_sva_31_2_mx0c1;
  wire GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c0;
  wire GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c1;
  wire GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c2;
  wire GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c4;
  wire GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c7;
  wire GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c9;
  wire GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c10;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c0;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c1;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c7;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c9;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx2;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c0;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c1;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c7;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c9;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx1;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c0;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c1;
  wire attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c0;
  wire attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c1;
  wire attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c5;
  wire attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c8;
  wire attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c10;
  wire GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c0;
  wire GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c1;
  wire GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c2;
  wire GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c3;
  wire GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c6;
  wire attention_abs_qr_35_0_lpi_1_dfm_mx0c1;
  wire [38:0] QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_dfm_1_38_0_1;
  wire RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c1;
  wire [2:0] TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3;
  wire [3:0] nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3;
  wire CACHE_UPDATE_LOOP_3_k_2_0_sva_1_mx0c1;
  wire GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c1;
  wire GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c2;
  wire [39:0] attention_abs_2_mux_2;
  wire [40:0] nl_attention_abs_2_mux_2;
  wire RMS_NORM_LOOP_2_and_29_ssc_1;
  wire RMS_NORM_LOOP_2_and_34_ssc_1;
  wire RMS_NORM_LOOP_2_2_and_32_ssc_mx0w3;
  wire RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_nor_1_ssc_1;
  wire RMS_NORM_LOOP_2_and_33_ssc_1;
  wire [38:0] QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_dfm_1_38_0_mx0w1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16_mx1;
  wire attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16_mx0c1;
  wire attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16_mx0c1;
  wire attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16_mx0c1;
  wire attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16_mx0c1;
  wire attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16_mx0c1;
  wire attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16_mx0c1;
  wire attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16_mx0c1;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c0;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c2;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c3;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c4;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c1;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c8;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1;
  wire attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c1;
  wire attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c6;
  wire attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0_mx0c1;
  wire [15:0] attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0_mx0w6;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16_mx0c1;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16_mx0c1;
  wire [23:0] LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48_mx0w2;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16_mx0w5;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16_mx1;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16_mx1;
  wire [2:0] LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_2;
  wire [3:0] nl_LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_2;
  wire [23:0] operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1;
  wire [24:0] nl_operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1;
  wire [23:0] operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1;
  wire [24:0] nl_operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1;
  wire [23:0] operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1;
  wire [24:0] nl_operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1;
  wire [23:0] RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1;
  wire GEMM_3D_FLOAT_LOOP_3_and_tmp_4_sva_mx0w2;
  wire GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_0_sva_mx0w3;
  wire GEMM_3D_FLOAT_LOOP_3_and_tmp_5_sva_mx0w2;
  wire GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_1_sva_mx0w3;
  wire GEMM_3D_FLOAT_LOOP_3_and_tmp_6_sva_mx0w1;
  wire GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva_mx0w3;
  wire GEMM_3D_FLOAT_LOOP_3_and_tmp_7_sva_mx0w1;
  wire GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva_mx0w3;
  wire [23:0] APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1;
  wire [23:0] APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1;
  wire [39:0] APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1;
  wire [40:0] nl_APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1;
  wire [39:0] APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1;
  wire [40:0] nl_APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1;
  wire [23:0] RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1;
  wire [15:0] RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c1;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c9;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx2;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx0c7;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx1;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx0c7;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx1;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c1;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c9;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx2;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx0c7;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx1;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx0c7;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx1;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx0c7;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx1;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c1;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c9;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx2;
  wire attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx0c7;
  wire [39:0] attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx1;
  wire [2:0] TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_15_sdt_1;
  wire [3:0] nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_15_sdt_1;
  wire GEMM_3D_FLOAT_LOOP_3_and_tmp_sva_mx0w0;
  wire GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva_mx0w0;
  wire GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva_mx0w0;
  wire GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva_mx0w0;
  wire GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva_mx0w0;
  wire GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva_mx0w0;
  wire GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva_mx0w0;
  wire GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva_mx0w0;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6_mx1;
  wire [38:0] SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1;
  wire [39:0] nl_SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1;
  wire [39:0] SF_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_psp_sva_1;
  wire [39:0] CM_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_ctmp_sva_1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9_mx1;
  wire [39:0] attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8_mx1;
  wire [39:0] SOFTMAX_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_cse_sva_1;
  wire [39:0] SOFTMAX_LOOP_4_acc_3_cse_sva_1;
  wire [40:0] nl_SOFTMAX_LOOP_4_acc_3_cse_sva_1;
  wire GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva_mx0w0;
  wire attention_abs_4_qr_35_0_lpi_1_dfm_mx0c1;
  wire [39:0] attention_abs_5_qr_sva_1;
  wire [40:0] nl_attention_abs_5_qr_sva_1;
  wire [39:0] attention_abs_6_mux_2;
  wire [40:0] nl_attention_abs_6_mux_2;
  wire RMS_NORM_LOOP_2_2_and_29_ssc_1;
  wire RMS_NORM_LOOP_2_2_and_34_ssc_1;
  wire RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_nor_1_ssc_1;
  wire RMS_NORM_LOOP_2_2_and_33_ssc_1;
  wire QUANTIZE_ACTIVATION_LOOP_3_1_nand_seb_1;
  wire [23:0] output_0_15_lpi_4_39_16_mx1;
  wire [23:0] output_0_0_lpi_4_39_16_mx1;
  wire [23:0] output_0_14_lpi_4_39_16_mx1;
  wire [23:0] output_0_1_lpi_4_39_16_mx1;
  wire [23:0] output_0_13_lpi_4_39_16_mx1;
  wire [23:0] output_0_2_lpi_4_39_16_mx1;
  wire [23:0] output_0_12_lpi_4_39_16_mx1;
  wire [23:0] output_0_3_lpi_4_39_16_mx1;
  wire [23:0] output_0_11_lpi_4_39_16_mx1;
  wire [23:0] output_0_4_lpi_4_39_16_mx1;
  wire [23:0] output_0_10_lpi_4_39_16_mx1;
  wire [23:0] output_0_5_lpi_4_39_16_mx1;
  wire [23:0] output_0_9_lpi_4_39_16_mx1;
  wire [23:0] output_0_6_lpi_4_39_16_mx1;
  wire [23:0] output_0_8_lpi_4_39_16_mx1;
  wire [23:0] output_0_7_lpi_4_39_16_mx1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_7_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_0_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_6_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_1_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_5_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_2_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_4_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_3_1;
  wire [23:0] operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1;
  wire [24:0] nl_operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1;
  reg [38:0] attention_abs_3_qr_sva_38_0;
  reg [38:0] attention_abs_5_qr_sva_38_0;
  reg [38:0] attention_abs_7_qr_sva_38_0;
  reg [13:0] output_0_7_sva_2_29_16;
  reg [13:0] output_0_8_sva_2_29_16;
  reg [13:0] output_0_6_sva_2_29_16;
  reg [13:0] output_0_9_sva_2_29_16;
  reg [13:0] output_0_5_sva_2_29_16;
  reg [13:0] output_0_10_sva_2_29_16;
  reg [13:0] output_0_4_sva_2_29_16;
  reg [13:0] output_0_11_sva_2_29_16;
  reg [13:0] output_0_3_sva_2_29_16;
  reg [13:0] output_0_12_sva_2_29_16;
  reg [13:0] output_0_2_sva_2_29_16;
  reg [13:0] output_0_13_sva_2_29_16;
  reg [13:0] output_0_1_sva_2_29_16;
  reg [13:0] output_0_14_sva_2_29_16;
  reg [13:0] output_0_0_sva_2_29_16;
  reg [13:0] output_0_15_sva_2_29_16;
  wire attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_39;
  wire [38:0] attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_38_0;
  reg attention_abs_qr_35_0_lpi_1_dfm_35;
  reg [34:0] attention_abs_qr_35_0_lpi_1_dfm_34_0;
  reg attention_abs_4_qr_35_0_lpi_1_dfm_35;
  reg [34:0] attention_abs_4_qr_35_0_lpi_1_dfm_34_0;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_15_8;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_15_8;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_15_8;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_15_8;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_15_8;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_15_8;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_8;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_15_8;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_15_8;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_15_8;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_15_8;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_15_8;
  wire [11:0] operator_40_24_true_AC_TRN_AC_WRAP_1_conc_1_itm_11_0;
  wire [8:0] operator_40_24_true_AC_TRN_AC_WRAP_1_conc_3_itm_8_0;
  wire RMS_NORM_LOOP_1_1_or_3_ssc;
  wire RMS_NORM_LOOP_1_1_or_1_ssc;
  reg reg_rms_norm_16_div_cmp_b_ftd_1;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd;
  reg [38:0] reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1;
  reg [2:0] reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd;
  reg [2:0] reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1;
  reg reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2;
  reg [7:0] reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3;
  wire attention_2_1_16_16_4_4_q_proj_and_4_ssc;
  reg reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd;
  reg reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_1;
  reg reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_2;
  reg reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_3;
  reg reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_4;
  reg reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_5;
  reg reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_6;
  reg reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_7;
  reg [7:0] reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd;
  reg [7:0] reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd;
  wire and_581_ssc;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_nand_seb;
  wire and_585_seb;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_1_ssc;
  reg LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4;
  reg [3:0] LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_2_or_1_cse;
  wire rms_norm_16_variance_or_1_cse;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_cse;
  wire attention_2_1_16_16_4_4_attn_output_and_14_cse;
  wire attention_2_1_16_16_4_4_attn_output_and_13_cse;
  wire attention_2_1_16_16_4_4_attn_output_and_16_cse;
  wire attention_2_1_16_16_4_4_attn_output_and_15_cse;
  wire attention_2_1_16_16_4_4_attn_output_and_18_cse;
  wire attention_2_1_16_16_4_4_attn_output_and_17_cse;
  wire attention_2_1_16_16_4_4_q_proj_re_and_cse;
  wire attention_2_1_16_16_4_4_k_proj_re_and_1_cse;
  wire nor_1053_cse;
  wire nor_1044_cse;
  wire nor_1045_cse;
  wire nor_1138_m1c;
  reg [7:0] LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_47_40;
  reg [7:0] reg_rms_norm_16_div_cmp_a_ftd_1_15_8;
  wire GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_8_seb;
  wire or_1667_ssc;
  wire attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_39;
  wire [38:0] attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_38_0;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_7;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_6;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_5;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_4;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_3;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_2;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_0;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_7;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_6;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_5;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_4;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_3;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_2;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_0;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_7;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_6;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_5;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_4;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_3;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_2;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_0;
  reg attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_39;
  reg [38:0] attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_38_0;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0;
  wire RMS_NORM_LOOP_1_1_or_2_ssc;
  wire nor_1314_cse;
  wire mux_1513_cse;
  wire CACHE_UPDATE_LOOP_3_or_cse;
  wire CACHE_UPDATE_LOOP_3_or_1_cse;
  wire RMS_NORM_LOOP_1_1_or_5_cse;
  wire compute_sqrt_for_i_and_2_cse;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_and_31_cse;
  wire [23:0] attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
  wire RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
  wire attention_2_1_16_16_4_4_quantized_hidden_states_and_3_ssc;
  reg attention_2_1_16_16_4_4_quantized_hidden_states_0_7_sva_7;
  wire attention_2_1_16_16_4_4_quantized_hidden_states_and_2_ssc;
  reg attention_2_1_16_16_4_4_quantized_hidden_states_0_8_sva_7;
  wire attention_2_1_16_16_4_4_quantized_hidden_states_and_1_ssc;
  reg attention_2_1_16_16_4_4_quantized_hidden_states_0_6_sva_7;
  wire attention_2_1_16_16_4_4_quantized_hidden_states_and_ssc;
  reg attention_2_1_16_16_4_4_quantized_hidden_states_0_9_sva_7;
  reg attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_15;
  reg [2:0] attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_14_12;
  reg [2:0] attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_11_9;
  reg attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_8;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0;
  wire [7:0] apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
  wire [7:0] apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
  wire [7:0] attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_15_8;
  wire attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_0;
  wire [7:0] attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_15_8;
  wire attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_0;
  wire [7:0] attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_15_8;
  wire attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_0;
  wire [7:0] attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_15_8;
  wire attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_0;
  wire [7:0] attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_15_8;
  wire attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_0;
  wire [7:0] attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_15_8;
  wire attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_0;
  wire [7:0] attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_15_8;
  wire attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_0;
  wire [7:0] attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_15_8;
  wire [7:0] attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_15_8;
  wire attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_0;
  wire [7:0] attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_15_8;
  wire attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_0;
  wire [7:0] attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_15_8;
  wire attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_0;
  wire [7:0] attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_15_8;
  wire attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_0;
  wire [7:0] attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_15_8;
  wire [7:0] attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_15_8;
  wire nor_1228_ssc;
  wire attention_2_1_16_16_4_4_q_proj_and_5_ssc;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_7;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_6;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_5;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_4;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_3;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_2;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_1;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_0;
  reg input_0_13_sva_1_39;
  reg [38:0] input_0_13_sva_1_38_0;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_7;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_6;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_5;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_4;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_3;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_2;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_1;
  reg attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_0;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_7;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_6;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_5;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_4;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_3;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_2;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_1;
  reg attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_0;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_7;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_6;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_5;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_4;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_3;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_2;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_1;
  reg attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_0;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_7;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_6;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_5;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_4;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_3;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_2;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_1;
  reg attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_0;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_7;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_6;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_5;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_4;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_3;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_2;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_1;
  reg attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_0;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_7;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_6;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_5;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_4;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_3;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_2;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_1;
  reg attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_0;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8;
  reg attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_7;
  reg attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_6;
  reg attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_5;
  reg attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_4;
  reg attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_3;
  reg attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_2;
  reg attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_1;
  reg attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_0;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_7;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_6;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_5;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_4;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_3;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_2;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_1;
  reg attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_0;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_7;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_6;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_5;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_4;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_3;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_2;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_1;
  reg attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_0;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_7;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_6;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_5;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_4;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_3;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_2;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_1;
  reg attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_0;
  reg [7:0] attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_7;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_6;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_5;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_4;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_3;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_2;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_1;
  reg attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_0;
  reg [7:0] attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_8;
  reg [7:0] attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_8;
  reg [7:0] apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_8;
  reg [7:0] apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_8;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_1_and_29_ssc;
  reg [7:0] LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8;
  wire attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_0;
  reg reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_cse;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_cse;
  wire RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
  wire and_474_rgt;
  wire and_476_rgt;
  wire and_480_rgt;
  wire for_for_and_14_rgt;
  wire for_for_and_15_rgt;
  wire for_for_and_16_rgt;
  wire for_for_and_17_rgt;
  wire and_485_rgt;
  wire and_486_rgt;
  wire for_for_or_1_rgt;
  wire and_745_ssc;
  reg input_0_13_sva_2_39;
  reg [38:0] input_0_13_sva_2_38_0;
  wire [7:0] apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
  wire attention_abs_qr_35_0_lpi_1_dfm_mx1_35;
  wire [33:0] attention_abs_qr_35_0_lpi_1_dfm_mx1_34_1;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_7;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_6;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_5;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_4;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_3;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_2;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_1;
  reg attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_0;
  wire and_303_ssc;
  wire compute_sqrt_guess_or_1_ssc;
  wire and_315_ssc;
  reg operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_34;
  reg [33:0] operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_33_0;
  wire QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_and_ssc;
  reg QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39;
  reg [38:0] QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0;
  wire compute_sqrt_guess_and_ssc;
  reg compute_sqrt_guess_sva_34;
  reg [33:0] compute_sqrt_guess_sva_33_0;
  reg [7:0] attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_15_8;
  reg [7:0] apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_8;
  wire compute_sqrt_1_guess_and_ssc;
  reg compute_sqrt_1_guess_sva_34;
  reg [33:0] compute_sqrt_1_guess_sva_33_0;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_or_11_cse;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_or_12_cse;
  wire attention_2_1_16_16_4_4_q_embed_and_25_cse;
  wire attention_2_1_16_16_4_4_q_embed_and_27_cse;
  wire attention_2_1_16_16_4_4_q_embed_and_29_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse;
  reg reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse;
  wire attention_2_1_16_16_4_4_k_proj_re_or_cse;
  wire attention_2_1_16_16_4_4_k_proj_re_or_17_cse;
  wire RMS_NORM_LOOP_2_2_i_and_9_cse;
  wire attention_2_1_16_16_4_4_k_proj_re_and_91_cse;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse;
  wire GEMM_3D_FLOAT_LOOP_4_l_or_2_cse;
  reg input_0_2_sva_1_39;
  reg [38:0] input_0_2_sva_1_38_0;
  wire [7:0] APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8;
  wire and_699_ssc;
  reg input_0_2_sva_2_39;
  reg [38:0] input_0_2_sva_2_38_0;
  reg [7:0] apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_15_8;
  reg [7:0] apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_15_8;
  reg [7:0] apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_15_8;
  wire [7:0] apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
  wire attention_2_1_16_16_4_4_v_proj_and_2_cse;
  wire attention_2_1_16_16_4_4_q_embed_and_26_cse;
  wire attention_2_1_16_16_4_4_q_embed_and_28_cse;
  wire attention_2_1_16_16_4_4_q_embed_and_30_cse;
  wire operator_40_24_true_AC_TRN_AC_WRAP_1_and_4_cse;
  wire attention_2_1_16_16_4_4_q_proj_re_and_29_cse;
  wire attention_2_1_16_16_4_4_k_proj_re_and_65_cse;
  wire attention_2_1_16_16_4_4_v_proj_re_and_95_cse;
  wire attention_2_1_16_16_4_4_v_proj_and_30_cse;
  wire attention_2_1_16_16_4_4_attn_weights_and_52_cse;
  reg [7:0] reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_ftd;
  wire and_1055_ssc;
  wire and_1059_ssc;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_and_30_ssc;
  reg [7:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8;
  reg [7:0] attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_15_8;
  reg [7:0] output_0_1_lpi_3_15_8;
  reg [7:0] output_0_1_sva_2_15_8;
  wire [7:0] attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_15_8;
  wire attention_2_1_16_16_4_4_q_proj_and_23_cse;
  reg [7:0] reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_ftd;
  reg [7:0] strm_out_rsci_idat_17_10;
  reg operator_80_48_true_AC_TRN_AC_WRAP_operator_80_48_true_AC_TRN_AC_WRAP_slc_SOFTMAX_LOOP_4_sqr_56_1_itm_slc;
  reg [7:0] reg_QUANTIZE_ACTIVATION_LOOP_3_quantized_value_slc_63_32_cse_slc;
  reg [15:0] reg_RMS_NORM_LOOP_1_1_slc_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_mul_55_16_cse_1_slc;
  wire nand_302_cse;
  wire [7:0] RESHAPE_2D_TO_3D_LOOP_3_1_mux_13_cse;
  wire attention_2_1_16_16_4_4_q_embed_and_23_cse;
  wire attention_2_1_16_16_4_4_q_embed_and_24_cse;
  wire ATTN_2D_LOOP_3_mux_16_itm;
  wire [38:0] ATTN_2D_LOOP_3_mux_17_itm;
  wire GEMM_3D_FLOAT_LOOP_4_1_nand_itm;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_5_itm;
  wire mux_1512_itm;
  wire and_1034_itm;
  wire mux_1966_itm;
  wire and_1037_itm;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  wire [7:0] APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm;
  wire mux_1079_itm;
  wire RMS_NORM_LOOP_1_1_or_4_itm;
  wire [39:0] compute_sqrt_1_for_acc_1_itm_40_1_1;
  wire [39:0] compute_sqrt_for_acc_1_itm_40_1_1;
  wire QUANTIZE_ACTIVATION_LOOP_2_acc_4_itm_40_1;
  wire QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1;
  wire [39:0] APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1;
  wire [39:0] APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1;
  wire QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_itm_40_1;
  wire QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1;
  wire CACHE_UPDATE_LOOP_2_1_acc_2_itm_2_1;
  wire attention_max_attn_fixed_t_1_acc_1_itm_40_1;
  wire CACHE_UPDATE_LOOP_2_acc_2_itm_2_1;
  wire SOFTMAX_LOOP_3_acc_3_itm_40_1;
  reg [7:0] reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_1;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_2;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_3;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_4;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_5;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_6;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_7;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_8;
  reg [7:0] reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_1;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_2;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_3;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_4;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_5;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_6;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_7;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_8;
  reg [7:0] reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_1;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_2;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_3;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_4;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_5;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_6;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_7;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_8;
  wire GEMM_3D_FLOAT_LOOP_4_1_and_ssc;
  reg reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd;
  reg [38:0] reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_ssc;
  reg reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd;
  reg reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  reg [1:0] reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_and_ssc;
  reg reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd;
  reg [1:0] reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1;
  reg reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  wire GEMM_3D_FLOAT_LOOP_1_i_and_ssc;
  reg reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd;
  reg reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  wire APPLY_ROTARY_POS_EMB_LOOP_1_i_and_ssc;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_k_and_ssc;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_and_18_ssc;
  reg [2:0] reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd;
  reg [12:0] reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1;
  reg reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd;
  reg reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1;
  reg reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2;
  reg reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3;
  reg reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4;
  reg reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5;
  reg reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6;
  reg reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_and_17_ssc;
  reg [7:0] apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_8;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_7;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_6;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_5;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_4;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_3;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_2;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_1;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_0;
  wire and_1042_ssc;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_and_16_ssc;
  reg [7:0] apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_15_8;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_7;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_6;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_5;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_4;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_3;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_2;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_1;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_0;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
  wire [7:0] apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
  wire RMS_NORM_LOOP_1_1_nor_seb;
  wire and_1062_ssc;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_and_19_ssc;
  reg [7:0] apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_15_8;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_7;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_6;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_5;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_4;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_3;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_2;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_1;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_0;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_7;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_6;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_5;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_4;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_3;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_2;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_1;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_0;
  reg [7:0] apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_8;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_7;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_6;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_5;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_4;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_3;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_2;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_1;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_0;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_7;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_6;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_5;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_4;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_3;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_2;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_1;
  reg apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_0;
  wire apply_rotary_pos_emb_1_4_4_rotated_q_and_37_cse;
  wire attention_2_1_16_16_4_4_attn_output_and_25_cse;
  wire input_and_28_cse;
  wire output_and_64_cse;
  wire and_339_ssc;
  reg SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_39;
  reg [38:0] SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_38_0;
  wire and_329_ssc;
  wire and_334_ssc;
  reg SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_55;
  reg [38:0] SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_54_16;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_0;
  reg [2:0] attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_15_13;
  reg [12:0] attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0;
  reg [7:0] attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_15_8;
  reg attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_7;
  reg attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_6;
  reg attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_5;
  reg attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_4;
  reg attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_3;
  reg attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_2;
  reg attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_1;
  reg attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_0;
  wire [7:0] attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_15_8;
  wire attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_0;
  wire [2:0] attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_15_13;
  wire [12:0] attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0;
  reg [21:0] reg_rms_norm_16_div_cmp_b_ftd_59_38;
  reg [37:0] reg_rms_norm_16_div_cmp_b_ftd_37_0;
  reg LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_39;
  reg LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_38;
  reg LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_37;
  reg LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_36;
  reg LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_35;
  reg LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_34;
  reg LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_33;
  reg LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_32;
  reg reg_rms_norm_16_div_cmp_a_ftd_1_7;
  reg reg_rms_norm_16_div_cmp_a_ftd_1_6;
  reg reg_rms_norm_16_div_cmp_a_ftd_1_5;
  reg reg_rms_norm_16_div_cmp_a_ftd_1_4;
  reg reg_rms_norm_16_div_cmp_a_ftd_1_3;
  reg reg_rms_norm_16_div_cmp_a_ftd_1_2;
  reg reg_rms_norm_16_div_cmp_a_ftd_1_1;
  reg reg_rms_norm_16_div_cmp_a_ftd_1_0;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
  wire attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_0;
  wire RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_7;
  wire RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_6;
  wire RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_5;
  wire RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_4;
  wire RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_3;
  wire RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_2;
  wire RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_1;
  wire RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_0;
  wire [2:0] apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_13;
  wire [4:0] apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_12_8;
  reg [7:0] attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_8;
  reg attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_7;
  reg attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_6;
  reg attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_5;
  reg attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_4;
  reg attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_3;
  reg attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_2;
  reg attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_1;
  reg attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_0;
  reg [2:0] attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_13;
  reg [12:0] attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0;
  reg attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_7;
  reg attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_6;
  reg attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_5;
  reg attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_4;
  reg attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_3;
  reg attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_2;
  reg attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_1;
  reg attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_0;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_7;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_6;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_5;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_4;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_3;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_2;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_1;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_0;
  reg attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_7;
  reg attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_6;
  reg attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_5;
  reg attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_4;
  reg attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_3;
  reg attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_2;
  reg attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_1;
  reg attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_0;
  reg [2:0] apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_13;
  reg [4:0] apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_12_8;
  wire GEMM_3D_FLOAT_LOOP_1_or_ssc;
  wire and_1908_cse;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1;
  reg reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_1;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_0;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
  wire attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_0;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_7;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_6;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_5;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_4;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_3;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_2;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_1;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_0;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_7;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_6;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_5;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_4;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_3;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_2;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_1;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_0;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_7;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_6;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_5;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_4;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_3;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_2;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_1;
  reg apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_0;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
  wire apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_1;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_2;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_3;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_4;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_5;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_6;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_7;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_1;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_2;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_3;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_4;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_5;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_6;
  reg reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_7;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_1;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_2;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_3;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_4;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_5;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_6;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_7;
  reg APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7;
  reg APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6;
  reg APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5;
  reg APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4;
  reg APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3;
  reg APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2;
  reg APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1;
  reg APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0;
  reg attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_7;
  reg attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_6;
  reg attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_5;
  reg attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_4;
  reg attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_3;
  reg attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_2;
  reg attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_1;
  reg attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_0;
  reg output_0_1_lpi_3_7;
  reg output_0_1_lpi_3_6;
  reg output_0_1_lpi_3_5;
  reg output_0_1_lpi_3_4;
  reg output_0_1_lpi_3_3;
  reg output_0_1_lpi_3_2;
  reg output_0_1_lpi_3_1;
  reg output_0_1_lpi_3_0;
  reg output_0_1_sva_2_7;
  reg output_0_1_sva_2_6;
  reg output_0_1_sva_2_5;
  reg output_0_1_sva_2_4;
  reg output_0_1_sva_2_3;
  reg output_0_1_sva_2_2;
  reg output_0_1_sva_2_1;
  reg output_0_1_sva_2_0;
  wire attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_7;
  wire attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_6;
  wire attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_5;
  wire attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_4;
  wire attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_3;
  wire attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_2;
  wire attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_1;
  wire attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_0;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_7_cse;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_8_cse;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_9_cse;
  wire compute_sqrt_for_i_and_cse;
  wire compute_sqrt_for_i_and_4_cse;
  wire compute_sqrt_for_i_and_5_cse;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_1;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_2;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_3;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_4;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_5;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_6;
  reg reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_7;
  reg strm_out_rsci_idat_9;
  reg strm_out_rsci_idat_8;
  reg strm_out_rsci_idat_7;
  reg strm_out_rsci_idat_6;
  reg strm_out_rsci_idat_5;
  reg strm_out_rsci_idat_4;
  reg strm_out_rsci_idat_3;
  reg strm_out_rsci_idat_2;
  wire [43:0] z_out_13_71_28;
  wire [39:0] acc_3_cse_40_1;
  wire [40:0] nl_acc_3_cse_40_1;

  wire mux_778_nl;
  wire mux_777_nl;
  wire mux_776_nl;
  wire mux_775_nl;
  wire and_1481_nl;
  wire mux_774_nl;
  wire or_1677_nl;
  wire mux_773_nl;
  wire or_1676_nl;
  wire attention_2_1_16_16_4_4_q_embed_and_31_nl;
  wire attention_2_1_16_16_4_4_q_embed_and_32_nl;
  wire mux_786_nl;
  wire mux_785_nl;
  wire mux_784_nl;
  wire mux_783_nl;
  wire mux_782_nl;
  wire mux_781_nl;
  wire nor_728_nl;
  wire mux_780_nl;
  wire mux_779_nl;
  wire and_1383_nl;
  wire and_1485_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_1_and_32_nl;
  wire GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_4_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_1_and_34_nl;
  wire GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_6_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_1_and_30_nl;
  wire GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_2_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_1_and_40_nl;
  wire GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_12_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_1_and_42_nl;
  wire GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_14_nl;
  wire and_259_nl;
  wire mux_789_nl;
  wire and_267_nl;
  wire mux_797_nl;
  wire mux_796_nl;
  wire mux_795_nl;
  wire mux_794_nl;
  wire mux_793_nl;
  wire or_1734_nl;
  wire mux_791_nl;
  wire nand_307_nl;
  wire mux_790_nl;
  wire nand_308_nl;
  wire nand_309_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_1_and_38_nl;
  wire GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_10_nl;
  wire mux_804_nl;
  wire mux_803_nl;
  wire mux_802_nl;
  wire mux_801_nl;
  wire and_274_nl;
  wire mux_800_nl;
  wire mux_799_nl;
  wire nor_271_nl;
  wire mux_815_nl;
  wire mux_814_nl;
  wire or_1775_nl;
  wire or_1774_nl;
  wire mux_813_nl;
  wire mux_812_nl;
  wire or_1771_nl;
  wire mux_811_nl;
  wire nand_41_nl;
  wire[7:0] operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_nl;
  wire not_4947_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_1_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_2_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_3_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_4_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_5_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_6_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_7_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_8_nl;
  wire mux_838_nl;
  wire mux_850_nl;
  wire mux_849_nl;
  wire or_1803_nl;
  wire mux_848_nl;
  wire mux_847_nl;
  wire mux_846_nl;
  wire or_1802_nl;
  wire mux_845_nl;
  wire or_1799_nl;
  wire mux_844_nl;
  wire mux_843_nl;
  wire mux_842_nl;
  wire or_1798_nl;
  wire mux_840_nl;
  wire or_1792_nl;
  wire mux_853_nl;
  wire nor_977_nl;
  wire and_1562_nl;
  wire mux_852_nl;
  wire and_1561_nl;
  wire rms_norm_16_mux1h_nl;
  wire[3:0] rms_norm_16_mux1h_9_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_1_not_1_nl;
  wire mux_854_nl;
  wire SOFTMAX_LOOP_5_mux_24_nl;
  wire[23:0] LINEAR_FORWARD_NO_MUL_LOOP_2_2_mux1h_2_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_2_not_nl;
  wire nor_979_nl;
  wire mux_855_nl;
  wire or_1812_nl;
  wire and_1564_nl;
  wire mux_861_nl;
  wire mux_860_nl;
  wire mux_859_nl;
  wire mux_862_nl;
  wire mux_864_nl;
  wire mux_863_nl;
  wire rms_norm_16_mux1h_10_nl;
  wire[23:0] rms_norm_16_mux1h_6_nl;
  wire rms_norm_16_not_nl;
  wire[7:0] rms_norm_16_mux1h_7_nl;
  wire rms_norm_16_not_1_nl;
  wire rms_norm_16_mux1h_11_nl;
  wire rms_norm_16_mux1h_13_nl;
  wire rms_norm_16_mux1h_14_nl;
  wire rms_norm_16_mux1h_15_nl;
  wire rms_norm_16_mux1h_16_nl;
  wire rms_norm_16_mux1h_17_nl;
  wire rms_norm_16_mux1h_18_nl;
  wire rms_norm_16_mux1h_19_nl;
  wire mux_874_nl;
  wire mux_873_nl;
  wire nor_907_nl;
  wire mux_872_nl;
  wire mux_871_nl;
  wire mux_870_nl;
  wire or_85_nl;
  wire mux_878_nl;
  wire mux_877_nl;
  wire mux_876_nl;
  wire nor_294_nl;
  wire mux_882_nl;
  wire mux_881_nl;
  wire mux_880_nl;
  wire or_1840_nl;
  wire mux_886_nl;
  wire mux_885_nl;
  wire mux_884_nl;
  wire nor_301_nl;
  wire mux_902_nl;
  wire mux_901_nl;
  wire or_1857_nl;
  wire mux_900_nl;
  wire mux_899_nl;
  wire mux_898_nl;
  wire mux_897_nl;
  wire nor_980_nl;
  wire nor_981_nl;
  wire or_1854_nl;
  wire mux_896_nl;
  wire or_1853_nl;
  wire mux_895_nl;
  wire mux_894_nl;
  wire and_380_nl;
  wire mux_893_nl;
  wire mux_892_nl;
  wire mux_891_nl;
  wire nand_316_nl;
  wire or_1849_nl;
  wire mux_890_nl;
  wire mux_889_nl;
  wire mux_888_nl;
  wire or_1847_nl;
  wire mux_887_nl;
  wire or_1846_nl;
  wire or_1845_nl;
  wire mux_905_nl;
  wire or_3156_nl;
  wire or_3157_nl;
  wire mux_948_nl;
  wire nor_985_nl;
  wire mux_947_nl;
  wire and_1566_nl;
  wire nor_986_nl;
  wire mux_946_nl;
  wire mux_945_nl;
  wire mux_944_nl;
  wire mux_943_nl;
  wire mux_942_nl;
  wire mux_941_nl;
  wire mux_940_nl;
  wire mux_939_nl;
  wire mux_938_nl;
  wire mux_935_nl;
  wire mux_934_nl;
  wire mux_933_nl;
  wire mux_932_nl;
  wire mux_931_nl;
  wire mux_930_nl;
  wire mux_929_nl;
  wire mux_928_nl;
  wire mux_926_nl;
  wire mux_925_nl;
  wire mux_924_nl;
  wire mux_923_nl;
  wire mux_920_nl;
  wire mux_918_nl;
  wire mux_917_nl;
  wire mux_914_nl;
  wire mux_913_nl;
  wire mux_912_nl;
  wire mux_911_nl;
  wire mux_907_nl;
  wire rms_norm_16_variance_mux1h_nl;
  wire GEMM_3D_FLOAT_LOOP_4_1_mux_17_nl;
  wire[38:0] rms_norm_16_variance_mux1h_1_nl;
  wire[38:0] GEMM_3D_FLOAT_LOOP_4_1_mux_24_nl;
  wire mux_952_nl;
  wire nor_990_nl;
  wire mux_951_nl;
  wire or_1890_nl;
  wire or_1889_nl;
  wire mux_950_nl;
  wire or_3158_nl;
  wire nand_318_nl;
  wire and_1568_nl;
  wire mux_949_nl;
  wire nor_988_nl;
  wire nor_989_nl;
  wire mux_985_nl;
  wire nand_47_nl;
  wire mux_2236_nl;
  wire or_3206_nl;
  wire or_3207_nl;
  wire mux_981_nl;
  wire or_3159_nl;
  wire mux_980_nl;
  wire mux_979_nl;
  wire mux_978_nl;
  wire or_1923_nl;
  wire or_1922_nl;
  wire or_1920_nl;
  wire mux_977_nl;
  wire or_1919_nl;
  wire or_1918_nl;
  wire or_3160_nl;
  wire mux_976_nl;
  wire or_1916_nl;
  wire nand_321_nl;
  wire mux_974_nl;
  wire mux_973_nl;
  wire mux_972_nl;
  wire mux_971_nl;
  wire mux_970_nl;
  wire mux_969_nl;
  wire nor_991_nl;
  wire mux_966_nl;
  wire mux_965_nl;
  wire mux_964_nl;
  wire mux_963_nl;
  wire mux_961_nl;
  wire nand_319_nl;
  wire mux_959_nl;
  wire mux_957_nl;
  wire or_1901_nl;
  wire or_1899_nl;
  wire nand_46_nl;
  wire mux_956_nl;
  wire mux_955_nl;
  wire mux_954_nl;
  wire or_1898_nl;
  wire or_1895_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_8_nl;
  wire[1:0] LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_9_nl;
  wire[1:0] QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_1_nl;
  wire[1:0] QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux_nl;
  wire and_1238_nl;
  wire nor_1322_nl;
  wire mux_2232_nl;
  wire mux_2231_nl;
  wire mux_2230_nl;
  wire and_426_nl;
  wire mux_984_nl;
  wire mux_983_nl;
  wire nor_996_nl;
  wire mux_982_nl;
  wire compute_sqrt_for_i_mux1h_nl;
  wire mux_2229_nl;
  wire mux_2228_nl;
  wire mux_2227_nl;
  wire nor_1311_nl;
  wire[1:0] compute_sqrt_for_i_nand_1_nl;
  wire[1:0] compute_sqrt_for_i_mux1h_1_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_not_2_nl;
  wire compute_sqrt_for_i_mux1h_2_nl;
  wire compute_sqrt_for_i_or_nl;
  wire[23:0] INIT_2D_MEM_LOOP_2_1_and_nl;
  wire[23:0] INIT_2D_MEM_LOOP_2_1_mux1h_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_37_nl;
  wire[22:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_69_nl;
  wire nor_1225_nl;
  wire mux_2081_nl;
  wire mux_2080_nl;
  wire nand_373_nl;
  wire mux_2079_nl;
  wire nor_576_nl;
  wire or_2777_nl;
  wire mux_2077_nl;
  wire or_2775_nl;
  wire and_1110_nl;
  wire and_1115_nl;
  wire nor_1323_nl;
  wire mux_2076_nl;
  wire nand_96_nl;
  wire mux_2075_nl;
  wire mux_2074_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_4_mux_17_nl;
  wire[39:0] SOFTMAX_LOOP_4_x_acc_2_nl;
  wire[40:0] nl_SOFTMAX_LOOP_4_x_acc_2_nl;
  wire[39:0] SOFTMAX_LOOP_4_x_mux_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_4_1_mux_18_nl;
  wire mux_1063_nl;
  wire mux_1062_nl;
  wire mux_1061_nl;
  wire mux_1060_nl;
  wire mux_1059_nl;
  wire mux_1058_nl;
  wire mux_1057_nl;
  wire mux_1056_nl;
  wire mux_1055_nl;
  wire mux_1054_nl;
  wire mux_1053_nl;
  wire mux_1050_nl;
  wire or_1996_nl;
  wire mux_1049_nl;
  wire mux_1048_nl;
  wire or_1994_nl;
  wire mux_1047_nl;
  wire mux_1046_nl;
  wire mux_1045_nl;
  wire mux_1043_nl;
  wire mux_1042_nl;
  wire mux_1072_nl;
  wire mux_1071_nl;
  wire mux_1070_nl;
  wire nand_328_nl;
  wire mux_1069_nl;
  wire mux_1068_nl;
  wire or_2016_nl;
  wire or_2015_nl;
  wire or_2014_nl;
  wire mux_1067_nl;
  wire mux_1066_nl;
  wire or_2013_nl;
  wire mux_1065_nl;
  wire or_2008_nl;
  wire mux_1064_nl;
  wire or_2007_nl;
  wire or_2006_nl;
  wire nand_329_nl;
  wire RMS_NORM_LOOP_2_mux_22_nl;
  wire QUANTIZE_ACTIVATION_LOOP_3_quantized_value_mux_nl;
  wire[38:0] RMS_NORM_LOOP_2_mux_24_nl;
  wire[38:0] QUANTIZE_ACTIVATION_LOOP_3_quantized_value_mux_1_nl;
  wire[39:0] for_for_mux1h_5_nl;
  wire for_for_for_for_nand_nl;
  wire for_for_and_24_nl;
  wire attention_2_1_16_16_4_4_attn_output_2D_not_nl;
  wire[39:0] for_for_mux1h_6_nl;
  wire attention_2_1_16_16_4_4_attn_output_2D_not_3_nl;
  wire mux_1099_nl;
  wire mux_1097_nl;
  wire mux_1095_nl;
  wire or_2048_nl;
  wire mux_1116_nl;
  wire mux_1115_nl;
  wire mux_1114_nl;
  wire GEMM_3D_FLOAT_LOOP_3_1_and_36_nl;
  wire[38:0] GEMM_3D_FLOAT_LOOP_3_1_and_52_nl;
  wire for_for_and_22_nl;
  wire mux_1119_nl;
  wire mux_1118_nl;
  wire mux_1117_nl;
  wire or_2081_nl;
  wire or_2080_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_1_and_28_nl;
  wire GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_nl;
  wire and_521_nl;
  wire and_523_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_1_and_29_nl;
  wire GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_1_nl;
  wire and_527_nl;
  wire and_529_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_1_and_31_nl;
  wire GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_3_nl;
  wire and_531_nl;
  wire and_533_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_1_and_33_nl;
  wire GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_5_nl;
  wire and_535_nl;
  wire and_537_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_1_and_35_nl;
  wire GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_7_nl;
  wire and_539_nl;
  wire and_541_nl;
  wire[39:0] mux_nl;
  wire[39:0] for_for_or_3_nl;
  wire[39:0] for_for_mux1h_13_nl;
  wire for_for_or_4_nl;
  wire for_for_and_28_nl;
  wire or_nl;
  wire nor_nl;
  wire mux_1133_nl;
  wire or_2087_nl;
  wire[39:0] mux1h_nl;
  wire or_3215_nl;
  wire not_4622_nl;
  wire[39:0] mux1h_1_nl;
  wire or_3216_nl;
  wire not_4624_nl;
  wire[39:0] mux1h_2_nl;
  wire or_3217_nl;
  wire not_4626_nl;
  wire mux_1211_nl;
  wire mux_1210_nl;
  wire mux_1209_nl;
  wire mux_1208_nl;
  wire mux_1212_nl;
  wire nor_1046_nl;
  wire and_1597_nl;
  wire mux_1235_nl;
  wire mux_1234_nl;
  wire mux_1233_nl;
  wire mux_1232_nl;
  wire mux_1231_nl;
  wire mux_1230_nl;
  wire mux_1228_nl;
  wire mux_1227_nl;
  wire mux_1226_nl;
  wire mux_1225_nl;
  wire mux_1224_nl;
  wire mux_1223_nl;
  wire or_2152_nl;
  wire or_2151_nl;
  wire or_2150_nl;
  wire mux_1222_nl;
  wire mux_1221_nl;
  wire mux_1220_nl;
  wire mux_1217_nl;
  wire mux_1216_nl;
  wire or_2145_nl;
  wire mux_1215_nl;
  wire mux_1214_nl;
  wire mux_1213_nl;
  wire or_2142_nl;
  wire or_2140_nl;
  wire or_2138_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_7_nl;
  wire[3:0] LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_4_nl;
  wire[3:0] LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_10_nl;
  wire mux_1310_nl;
  wire attention_2_1_16_16_4_4_q_proj_attention_2_1_16_16_4_4_q_proj_mux_12_nl;
  wire mux_1308_nl;
  wire or_3174_nl;
  wire nand_344_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_1_and_2_nl;
  wire[2:0] RMS_NORM_LOOP_2_2_i_mux1h_3_nl;
  wire RMS_NORM_LOOP_2_2_i_not_2_nl;
  wire RMS_NORM_LOOP_2_2_i_mux1h_6_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_and_10_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_nl;
  wire INIT_2D_MEM_LOOP_2_mux_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_38_nl;
  wire INIT_2D_MEM_LOOP_2_mux_10_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_39_nl;
  wire INIT_2D_MEM_LOOP_2_mux_11_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_40_nl;
  wire INIT_2D_MEM_LOOP_2_mux_12_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_41_nl;
  wire INIT_2D_MEM_LOOP_2_mux_13_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_42_nl;
  wire INIT_2D_MEM_LOOP_2_mux_14_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_43_nl;
  wire INIT_2D_MEM_LOOP_2_mux_15_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_44_nl;
  wire INIT_2D_MEM_LOOP_2_mux_16_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_1_nl;
  wire INIT_2D_MEM_LOOP_2_mux_1_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_24_nl;
  wire INIT_2D_MEM_LOOP_2_mux_17_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_nl;
  wire INIT_2D_MEM_LOOP_2_mux_18_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_26_nl;
  wire INIT_2D_MEM_LOOP_2_mux_19_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_27_nl;
  wire INIT_2D_MEM_LOOP_2_mux_20_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_28_nl;
  wire INIT_2D_MEM_LOOP_2_mux_21_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_29_nl;
  wire INIT_2D_MEM_LOOP_2_mux_22_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_30_nl;
  wire INIT_2D_MEM_LOOP_2_mux_23_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_2_nl;
  wire INIT_2D_MEM_LOOP_2_mux_2_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_10_nl;
  wire INIT_2D_MEM_LOOP_2_mux_24_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_11_nl;
  wire INIT_2D_MEM_LOOP_2_mux_25_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_12_nl;
  wire INIT_2D_MEM_LOOP_2_mux_26_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_13_nl;
  wire INIT_2D_MEM_LOOP_2_mux_27_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_14_nl;
  wire INIT_2D_MEM_LOOP_2_mux_28_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_15_nl;
  wire INIT_2D_MEM_LOOP_2_mux_29_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_16_nl;
  wire INIT_2D_MEM_LOOP_2_mux_30_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_3_nl;
  wire INIT_2D_MEM_LOOP_2_mux_3_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_17_nl;
  wire INIT_2D_MEM_LOOP_2_mux_31_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_18_nl;
  wire INIT_2D_MEM_LOOP_2_mux_32_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_19_nl;
  wire INIT_2D_MEM_LOOP_2_mux_33_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_20_nl;
  wire INIT_2D_MEM_LOOP_2_mux_34_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_21_nl;
  wire INIT_2D_MEM_LOOP_2_mux_35_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_22_nl;
  wire INIT_2D_MEM_LOOP_2_mux_36_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_23_nl;
  wire INIT_2D_MEM_LOOP_2_mux_37_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_4_nl;
  wire INIT_2D_MEM_LOOP_2_mux_4_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_31_nl;
  wire INIT_2D_MEM_LOOP_2_mux_38_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_32_nl;
  wire INIT_2D_MEM_LOOP_2_mux_39_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_33_nl;
  wire INIT_2D_MEM_LOOP_2_mux_40_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_34_nl;
  wire INIT_2D_MEM_LOOP_2_mux_41_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_35_nl;
  wire INIT_2D_MEM_LOOP_2_mux_42_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_36_nl;
  wire INIT_2D_MEM_LOOP_2_mux_43_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_37_nl;
  wire INIT_2D_MEM_LOOP_2_mux_44_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_5_nl;
  wire INIT_2D_MEM_LOOP_2_mux_5_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_45_nl;
  wire INIT_2D_MEM_LOOP_2_mux_45_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_46_nl;
  wire INIT_2D_MEM_LOOP_2_mux_46_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_47_nl;
  wire INIT_2D_MEM_LOOP_2_mux_47_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_48_nl;
  wire INIT_2D_MEM_LOOP_2_mux_48_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_49_nl;
  wire INIT_2D_MEM_LOOP_2_mux_49_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_50_nl;
  wire INIT_2D_MEM_LOOP_2_mux_50_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_51_nl;
  wire INIT_2D_MEM_LOOP_2_mux_51_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_6_nl;
  wire INIT_2D_MEM_LOOP_2_mux_6_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_52_nl;
  wire INIT_2D_MEM_LOOP_2_mux_52_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_53_nl;
  wire INIT_2D_MEM_LOOP_2_mux_53_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_54_nl;
  wire INIT_2D_MEM_LOOP_2_mux_54_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_55_nl;
  wire INIT_2D_MEM_LOOP_2_mux_55_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_56_nl;
  wire INIT_2D_MEM_LOOP_2_mux_56_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_57_nl;
  wire INIT_2D_MEM_LOOP_2_mux_57_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_58_nl;
  wire INIT_2D_MEM_LOOP_2_mux_58_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_7_nl;
  wire INIT_2D_MEM_LOOP_2_mux_7_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_59_nl;
  wire INIT_2D_MEM_LOOP_2_mux_59_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_60_nl;
  wire INIT_2D_MEM_LOOP_2_mux_60_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_61_nl;
  wire INIT_2D_MEM_LOOP_2_mux_61_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_62_nl;
  wire INIT_2D_MEM_LOOP_2_mux_62_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_63_nl;
  wire INIT_2D_MEM_LOOP_2_mux_63_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_64_nl;
  wire INIT_2D_MEM_LOOP_2_mux_64_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_65_nl;
  wire INIT_2D_MEM_LOOP_2_mux_65_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_8_nl;
  wire INIT_2D_MEM_LOOP_2_mux_8_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_66_nl;
  wire INIT_2D_MEM_LOOP_2_mux_66_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_67_nl;
  wire INIT_2D_MEM_LOOP_2_mux_67_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_68_nl;
  wire INIT_2D_MEM_LOOP_2_mux_68_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_69_nl;
  wire INIT_2D_MEM_LOOP_2_mux_69_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_70_nl;
  wire INIT_2D_MEM_LOOP_2_mux_70_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_71_nl;
  wire INIT_2D_MEM_LOOP_2_mux_71_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_72_nl;
  wire INIT_2D_MEM_LOOP_2_mux_72_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_9_nl;
  wire INIT_2D_MEM_LOOP_2_mux_9_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_73_nl;
  wire INIT_2D_MEM_LOOP_2_mux_73_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_74_nl;
  wire INIT_2D_MEM_LOOP_2_mux_74_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_75_nl;
  wire INIT_2D_MEM_LOOP_2_mux_75_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_76_nl;
  wire INIT_2D_MEM_LOOP_2_mux_76_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_77_nl;
  wire INIT_2D_MEM_LOOP_2_mux_77_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_78_nl;
  wire INIT_2D_MEM_LOOP_2_mux_78_nl;
  wire INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_79_nl;
  wire INIT_2D_MEM_LOOP_2_mux_79_nl;
  wire mux_1434_nl;
  wire mux_1433_nl;
  wire or_2335_nl;
  wire mux_1432_nl;
  wire mux_1431_nl;
  wire mux_1430_nl;
  wire mux_1429_nl;
  wire mux_1428_nl;
  wire nor_1105_nl;
  wire or_2331_nl;
  wire mux_1638_nl;
  wire nand_71_nl;
  wire or_2563_nl;
  wire mux_1637_nl;
  wire mux_1636_nl;
  wire mux_1453_nl;
  wire mux_1452_nl;
  wire and_679_nl;
  wire QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_3_nl;
  wire QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_nl;
  wire RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_and_nl;
  wire QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_4_nl;
  wire QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_3_nl;
  wire CACHE_UPDATE_LOOP_3_k_and_1_nl;
  wire mux_1441_nl;
  wire nor_1109_nl;
  wire nor_1110_nl;
  wire mux_1457_nl;
  wire nor_1115_nl;
  wire mux_1456_nl;
  wire nand_350_nl;
  wire or_2355_nl;
  wire mux_1455_nl;
  wire nor_1116_nl;
  wire nor_1117_nl;
  wire mux_1454_nl;
  wire nor_1114_nl;
  wire GEMM_3D_FLOAT_LOOP_1_i_mux_1_nl;
  wire RMS_NORM_LOOP_2_2_and_36_nl;
  wire RMS_NORM_LOOP_2_2_mux1h_nl;
  wire or_594_nl;
  wire mux_1439_nl;
  wire or_2342_nl;
  wire mux_1438_nl;
  wire nand_348_nl;
  wire or_2341_nl;
  wire mux_1437_nl;
  wire or_2340_nl;
  wire or_2339_nl;
  wire mux_1490_nl;
  wire nand_126_nl;
  wire and_688_nl;
  wire and_693_nl;
  wire and_704_nl;
  wire and_709_nl;
  wire and_713_nl;
  wire and_717_nl;
  wire and_721_nl;
  wire and_725_nl;
  wire and_729_nl;
  wire and_733_nl;
  wire and_737_nl;
  wire and_741_nl;
  wire and_749_nl;
  wire and_753_nl;
  wire or_2443_nl;
  wire mux_1498_nl;
  wire mux_1497_nl;
  wire or_2429_nl;
  wire mux_1496_nl;
  wire or_2426_nl;
  wire mux_1495_nl;
  wire mux_1494_nl;
  wire mux_1493_nl;
  wire mux_1492_nl;
  wire nand_354_nl;
  wire nand_355_nl;
  wire mux_1511_nl;
  wire mux_1510_nl;
  wire or_2442_nl;
  wire mux_1509_nl;
  wire mux_1508_nl;
  wire mux_1507_nl;
  wire or_2441_nl;
  wire mux_1505_nl;
  wire or_2438_nl;
  wire nand_64_nl;
  wire mux_1504_nl;
  wire mux_1503_nl;
  wire or_2436_nl;
  wire nand_63_nl;
  wire mux_1502_nl;
  wire mux_1501_nl;
  wire mux_1500_nl;
  wire or_2431_nl;
  wire mux_1533_nl;
  wire mux_1532_nl;
  wire mux_1531_nl;
  wire mux_1530_nl;
  wire mux_1529_nl;
  wire or_2459_nl;
  wire mux_1528_nl;
  wire mux_1527_nl;
  wire or_2458_nl;
  wire mux_1526_nl;
  wire mux_1525_nl;
  wire mux_1524_nl;
  wire mux_1523_nl;
  wire mux_1521_nl;
  wire mux_1520_nl;
  wire mux_1518_nl;
  wire mux_1517_nl;
  wire or_2448_nl;
  wire or_2446_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_1_i_mux1h_5_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_2_and_1_nl;
  wire and_755_nl;
  wire nor_1136_nl;
  wire mux_1491_nl;
  wire nand_353_nl;
  wire and_757_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_1_i_or_nl;
  wire mux_1516_nl;
  wire nand_356_nl;
  wire mux_1515_nl;
  wire mux_1514_nl;
  wire mux_1537_nl;
  wire mux_1536_nl;
  wire nor_1141_nl;
  wire nor_1142_nl;
  wire nor_1143_nl;
  wire mux_1534_nl;
  wire or_2463_nl;
  wire or_2461_nl;
  wire mux_1541_nl;
  wire mux_1540_nl;
  wire mux_1539_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_4_nl;
  wire not_4557_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_8_nl;
  wire not_4558_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_12_nl;
  wire not_4559_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_16_nl;
  wire not_4560_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_20_nl;
  wire not_4561_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_21_nl;
  wire not_4562_nl;
  wire mux_1554_nl;
  wire and_1652_nl;
  wire mux_1552_nl;
  wire mux_1550_nl;
  wire or_2479_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_5_nl;
  wire and_779_nl;
  wire mux_1561_nl;
  wire mux_1560_nl;
  wire mux_1558_nl;
  wire mux_1556_nl;
  wire and_1653_nl;
  wire and_783_nl;
  wire and_790_nl;
  wire not_4472_nl;
  wire mux_1564_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_35_nl;
  wire not_4441_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_34_nl;
  wire not_4440_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_33_nl;
  wire not_4439_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_32_nl;
  wire not_4438_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_31_nl;
  wire not_4437_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_30_nl;
  wire not_4436_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_29_nl;
  wire not_4435_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_28_nl;
  wire not_4434_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_27_nl;
  wire not_4433_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_26_nl;
  wire not_4432_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_25_nl;
  wire not_4431_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_24_nl;
  wire not_4430_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_23_nl;
  wire not_4429_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_22_nl;
  wire not_4428_nl;
  wire mux_1581_nl;
  wire or_2494_nl;
  wire mux_1580_nl;
  wire or_2493_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_21_nl;
  wire not_4427_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_20_nl;
  wire not_4426_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_19_nl;
  wire not_4425_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_18_nl;
  wire not_4424_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_40_nl;
  wire not_4423_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_17_nl;
  wire not_4422_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_42_nl;
  wire not_4421_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_43_nl;
  wire not_4420_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_44_nl;
  wire not_4419_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_45_nl;
  wire not_4418_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_46_nl;
  wire not_4417_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_47_nl;
  wire not_4416_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_16_nl;
  wire not_4415_nl;
  wire GEMM_3D_FLOAT_LOOP_4_l_GEMM_3D_FLOAT_LOOP_4_l_mux_nl;
  wire GEMM_3D_FLOAT_LOOP_4_l_mux1h_13_nl;
  wire RMS_NORM_LOOP_1_1_or_nl;
  wire RMS_NORM_LOOP_1_1_mux1h_nl;
  wire RMS_NORM_LOOP_2_2_mux_23_nl;
  wire and_1254_nl;
  wire mux_2245_nl;
  wire mux_2244_nl;
  wire mux_2243_nl;
  wire mux_2242_nl;
  wire and_1810_nl;
  wire mux_2241_nl;
  wire nor_1320_nl;
  wire mux_2240_nl;
  wire nor_1316_nl;
  wire mux_2239_nl;
  wire and_1809_nl;
  wire nor_1321_nl;
  wire mux_2238_nl;
  wire or_3033_nl;
  wire or_3032_nl;
  wire GEMM_3D_FLOAT_LOOP_4_l_or_1_nl;
  wire or_2566_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_26_nl;
  wire and_939_nl;
  wire not_4471_nl;
  wire mux_1641_nl;
  wire or_3192_nl;
  wire mux_1640_nl;
  wire or_3191_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_28_nl;
  wire and_941_nl;
  wire not_4470_nl;
  wire mux_1644_nl;
  wire or_3195_nl;
  wire mux_1643_nl;
  wire or_3194_nl;
  wire or_2576_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_30_nl;
  wire and_943_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_nand_nl;
  wire mux_1660_nl;
  wire mux_1659_nl;
  wire mux_1657_nl;
  wire mux_1655_nl;
  wire nor_466_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_and_81_nl;
  wire and_945_nl;
  wire not_4469_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_32_nl;
  wire and_946_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_nand_2_nl;
  wire mux_1676_nl;
  wire mux_1675_nl;
  wire mux_1673_nl;
  wire mux_1671_nl;
  wire and_1684_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_and_83_nl;
  wire and_948_nl;
  wire not_4468_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_34_nl;
  wire and_949_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_nand_4_nl;
  wire mux_1692_nl;
  wire mux_1691_nl;
  wire mux_1689_nl;
  wire mux_1687_nl;
  wire or_2589_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_and_85_nl;
  wire and_951_nl;
  wire not_4467_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_36_nl;
  wire and_952_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_nand_6_nl;
  wire mux_1708_nl;
  wire mux_1707_nl;
  wire mux_1705_nl;
  wire mux_1703_nl;
  wire nand_367_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_and_87_nl;
  wire and_954_nl;
  wire not_4466_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_38_nl;
  wire and_955_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_nand_8_nl;
  wire mux_1724_nl;
  wire mux_1723_nl;
  wire mux_1721_nl;
  wire mux_1719_nl;
  wire and_1697_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_and_89_nl;
  wire and_957_nl;
  wire not_4465_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_40_nl;
  wire and_958_nl;
  wire not_4464_nl;
  wire mux_1727_nl;
  wire or_3197_nl;
  wire mux_1726_nl;
  wire nand_81_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_42_nl;
  wire and_960_nl;
  wire mux_1743_nl;
  wire mux_1742_nl;
  wire mux_1740_nl;
  wire mux_1738_nl;
  wire or_2611_nl;
  wire and_962_nl;
  wire not_4463_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_44_nl;
  wire and_963_nl;
  wire mux_1759_nl;
  wire mux_1758_nl;
  wire mux_1756_nl;
  wire mux_1754_nl;
  wire or_2617_nl;
  wire and_965_nl;
  wire not_4462_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_46_nl;
  wire and_966_nl;
  wire mux_1775_nl;
  wire mux_1774_nl;
  wire mux_1772_nl;
  wire mux_1770_nl;
  wire nor_500_nl;
  wire and_968_nl;
  wire not_4461_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_48_nl;
  wire and_969_nl;
  wire mux_1791_nl;
  wire mux_1790_nl;
  wire mux_1788_nl;
  wire mux_1786_nl;
  wire or_2492_nl;
  wire and_971_nl;
  wire not_4460_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_50_nl;
  wire and_972_nl;
  wire mux_1807_nl;
  wire mux_1806_nl;
  wire mux_1804_nl;
  wire mux_1802_nl;
  wire or_2497_nl;
  wire and_974_nl;
  wire not_4459_nl;
  wire mux_1811_nl;
  wire mux_1810_nl;
  wire or_2638_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_43_nl;
  wire not_4458_nl;
  wire mux_1816_nl;
  wire mux_1815_nl;
  wire mux_1814_nl;
  wire mux_1813_nl;
  wire or_2491_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_42_nl;
  wire not_4457_nl;
  wire mux_1825_nl;
  wire mux_1824_nl;
  wire mux_1823_nl;
  wire mux_1822_nl;
  wire or_2490_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_41_nl;
  wire not_4456_nl;
  wire mux_1834_nl;
  wire mux_1833_nl;
  wire mux_1832_nl;
  wire mux_1831_nl;
  wire nor_514_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_40_nl;
  wire not_4455_nl;
  wire mux_1843_nl;
  wire mux_1842_nl;
  wire mux_1841_nl;
  wire mux_1840_nl;
  wire and_1727_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_39_nl;
  wire not_4454_nl;
  wire mux_1852_nl;
  wire mux_1851_nl;
  wire mux_1850_nl;
  wire mux_1849_nl;
  wire or_2653_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_38_nl;
  wire not_4453_nl;
  wire mux_1861_nl;
  wire mux_1860_nl;
  wire mux_1859_nl;
  wire mux_1858_nl;
  wire nand_369_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_37_nl;
  wire not_4452_nl;
  wire mux_1870_nl;
  wire mux_1869_nl;
  wire mux_1868_nl;
  wire mux_1867_nl;
  wire and_1658_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_36_nl;
  wire not_4451_nl;
  wire mux_1878_nl;
  wire mux_1877_nl;
  wire mux_1876_nl;
  wire mux_1875_nl;
  wire mux_1874_nl;
  wire and_1733_nl;
  wire mux_1873_nl;
  wire or_2664_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_35_nl;
  wire not_4450_nl;
  wire mux_1887_nl;
  wire mux_1886_nl;
  wire mux_1885_nl;
  wire mux_1884_nl;
  wire nor_524_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_34_nl;
  wire not_4449_nl;
  wire mux_1896_nl;
  wire mux_1895_nl;
  wire mux_1894_nl;
  wire mux_1893_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_33_nl;
  wire not_4448_nl;
  wire mux_1905_nl;
  wire mux_1904_nl;
  wire mux_1903_nl;
  wire mux_1902_nl;
  wire or_2675_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_32_nl;
  wire not_4447_nl;
  wire mux_1914_nl;
  wire mux_1913_nl;
  wire mux_1912_nl;
  wire mux_1911_nl;
  wire nor_441_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_31_nl;
  wire not_4446_nl;
  wire mux_1923_nl;
  wire mux_1922_nl;
  wire mux_1921_nl;
  wire mux_1920_nl;
  wire and_1656_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_30_nl;
  wire not_4445_nl;
  wire mux_1932_nl;
  wire mux_1931_nl;
  wire mux_1930_nl;
  wire mux_1929_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_29_nl;
  wire not_4444_nl;
  wire mux_1941_nl;
  wire mux_1940_nl;
  wire mux_1939_nl;
  wire mux_1938_nl;
  wire or_2487_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_66_nl;
  wire and_1025_nl;
  wire not_4563_nl;
  wire mux_1946_nl;
  wire nor_533_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_67_nl;
  wire and_1031_nl;
  wire not_4564_nl;
  wire mux_1947_nl;
  wire nor_535_nl;
  wire mux_1965_nl;
  wire mux_1964_nl;
  wire mux_1962_nl;
  wire mux_1961_nl;
  wire mux_1960_nl;
  wire mux_1959_nl;
  wire mux_1958_nl;
  wire mux_1957_nl;
  wire mux_1954_nl;
  wire nor_540_nl;
  wire mux_1950_nl;
  wire or_2696_nl;
  wire mux_1949_nl;
  wire mux_1948_nl;
  wire or_2695_nl;
  wire[7:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_68_nl;
  wire[7:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_118_nl;
  wire not_4443_nl;
  wire[7:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_69_nl;
  wire[7:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_119_nl;
  wire not_4565_nl;
  wire mux_1973_nl;
  wire mux_1972_nl;
  wire and_1753_nl;
  wire mux_1971_nl;
  wire mux_1970_nl;
  wire nor_1203_nl;
  wire nor_1204_nl;
  wire and_1749_nl;
  wire mux_1969_nl;
  wire nor_1201_nl;
  wire nor_1202_nl;
  wire nor_1206_nl;
  wire mux_1968_nl;
  wire mux_1967_nl;
  wire and_1754_nl;
  wire nor_1208_nl;
  wire mux_1985_nl;
  wire mux_1984_nl;
  wire mux_1983_nl;
  wire mux_1982_nl;
  wire nor_551_nl;
  wire mux_1978_nl;
  wire mux_1977_nl;
  wire mux_1976_nl;
  wire or_2712_nl;
  wire mux_1975_nl;
  wire[7:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_70_nl;
  wire not_5074_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_128_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_129_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_130_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_131_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_132_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_133_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_134_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_135_nl;
  wire mux_1998_nl;
  wire mux_1997_nl;
  wire mux_1996_nl;
  wire mux_1995_nl;
  wire mux_1994_nl;
  wire nor_552_nl;
  wire mux_1992_nl;
  wire mux_1991_nl;
  wire mux_1989_nl;
  wire mux_1988_nl;
  wire or_2716_nl;
  wire mux_1987_nl;
  wire or_2715_nl;
  wire[7:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_71_nl;
  wire not_5066_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_120_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_121_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_122_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_123_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_124_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_125_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_126_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_127_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_72_nl;
  wire not_4566_nl;
  wire mux_2012_nl;
  wire mux_2011_nl;
  wire nand_93_nl;
  wire mux_2010_nl;
  wire mux_2009_nl;
  wire mux_2008_nl;
  wire mux_2007_nl;
  wire nand_92_nl;
  wire mux_2006_nl;
  wire mux_2005_nl;
  wire mux_2003_nl;
  wire mux_2002_nl;
  wire and_1759_nl;
  wire mux_2001_nl;
  wire mux_2000_nl;
  wire or_2720_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_73_nl;
  wire not_4567_nl;
  wire mux_2022_nl;
  wire mux_2021_nl;
  wire mux_2020_nl;
  wire mux_2019_nl;
  wire mux_2018_nl;
  wire or_2733_nl;
  wire and_1763_nl;
  wire mux_2017_nl;
  wire mux_2016_nl;
  wire mux_2033_nl;
  wire mux_2031_nl;
  wire mux_2030_nl;
  wire mux_2029_nl;
  wire mux_2028_nl;
  wire or_2741_nl;
  wire mux_2027_nl;
  wire[7:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_74_nl;
  wire[7:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_nl;
  wire not_5054_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_117_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_67_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_152_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_88_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_153_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_89_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_154_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_90_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_155_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_91_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_156_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_92_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_157_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_93_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_158_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_94_nl;
  wire mux_2036_nl;
  wire nor_410_nl;
  wire[2:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_75_nl;
  wire not_4569_nl;
  wire[4:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_116_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_144_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_145_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_146_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_147_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_148_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_149_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_150_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_151_nl;
  wire not_5062_nl;
  wire mux_2037_nl;
  wire and_1626_nl;
  wire[7:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_76_nl;
  wire not_5088_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_136_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_137_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_138_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_139_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_140_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_141_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_142_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux1h_143_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_77_nl;
  wire and_1064_nl;
  wire not_4571_nl;
  wire mux_2038_nl;
  wire nor_796_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_78_nl;
  wire and_1066_nl;
  wire not_4572_nl;
  wire mux_2039_nl;
  wire and_1420_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_79_nl;
  wire and_1068_nl;
  wire not_4573_nl;
  wire mux_2040_nl;
  wire and_1613_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_80_nl;
  wire and_1071_nl;
  wire and_1074_nl;
  wire not_4574_nl;
  wire mux_2051_nl;
  wire mux_2049_nl;
  wire mux_2048_nl;
  wire mux_2047_nl;
  wire mux_2046_nl;
  wire or_2751_nl;
  wire mux_2045_nl;
  wire and_1660_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_81_nl;
  wire and_1075_nl;
  wire not_4575_nl;
  wire mux_2052_nl;
  wire or_2753_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_82_nl;
  wire and_1081_nl;
  wire not_4576_nl;
  wire mux_2053_nl;
  wire or_2281_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_83_nl;
  wire and_1083_nl;
  wire not_4577_nl;
  wire mux_2054_nl;
  wire or_2292_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux1h_84_nl;
  wire and_1086_nl;
  wire not_4578_nl;
  wire mux_2055_nl;
  wire or_2756_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_51_nl;
  wire and_1089_nl;
  wire mux_2056_nl;
  wire or_2757_nl;
  wire not_4414_nl;
  wire mux_2059_nl;
  wire or_3200_nl;
  wire mux_2058_nl;
  wire and_1090_nl;
  wire mux_2057_nl;
  wire nor_1217_nl;
  wire or_3201_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_52_nl;
  wire not_4413_nl;
  wire mux_2063_nl;
  wire or_2764_nl;
  wire mux_2062_nl;
  wire or_2763_nl;
  wire mux_2061_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_53_nl;
  wire and_1097_nl;
  wire mux_2064_nl;
  wire or_2765_nl;
  wire not_4412_nl;
  wire mux_2068_nl;
  wire mux_2065_nl;
  wire nand_370_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_54_nl;
  wire not_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_55_nl;
  wire not_4579_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_56_nl;
  wire[23:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_36_nl;
  wire not_4580_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_57_nl;
  wire[23:0] LINEAR_FORWARD_NO_MUL_LOOP_2_mux_33_nl;
  wire[23:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_38_nl;
  wire not_4581_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_58_nl;
  wire[23:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_39_nl;
  wire not_4582_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_59_nl;
  wire not_4583_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_60_nl;
  wire not_4584_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_61_nl;
  wire not_4585_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_62_nl;
  wire not_4586_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_63_nl;
  wire not_4587_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux1h_64_nl;
  wire not_4588_nl;
  wire mux_2088_nl;
  wire mux_2087_nl;
  wire mux_2086_nl;
  wire mux_1542_nl;
  wire nand_357_nl;
  wire QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_nl;
  wire mux_2099_nl;
  wire mux_2098_nl;
  wire or_2799_nl;
  wire mux_2097_nl;
  wire mux_2096_nl;
  wire mux_2095_nl;
  wire mux_2094_nl;
  wire mux_2093_nl;
  wire mux_2091_nl;
  wire mux_2090_nl;
  wire or_2787_nl;
  wire or_2786_nl;
  wire QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_1_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_APPLY_ROTARY_POS_EMB_LOOP_3_nor_nl;
  wire QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_or_2_nl;
  wire[7:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_66_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_74_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_75_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_76_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_77_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_78_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_79_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_80_nl;
  wire[7:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_61_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_81_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_82_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_83_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_84_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_85_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_86_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_87_nl;
  wire mux_2102_nl;
  wire nand_283_nl;
  wire mux_2104_nl;
  wire mux_2103_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_32_nl;
  wire[2:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_70_nl;
  wire[2:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_71_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_72_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_50_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_51_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_52_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_53_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_54_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_55_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_56_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_57_nl;
  wire mux_2108_nl;
  wire nand_285_nl;
  wire or_3153_nl;
  wire mux_2107_nl;
  wire or_2828_nl;
  wire and_1184_nl;
  wire mux_2109_nl;
  wire GEMM_3D_FLOAT_LOOP_3_1_mux_4_nl;
  wire mux_2127_nl;
  wire mux_2126_nl;
  wire mux_2125_nl;
  wire mux_2124_nl;
  wire mux_2123_nl;
  wire mux_2122_nl;
  wire mux_2120_nl;
  wire mux_2114_nl;
  wire or_2840_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_and_7_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_and_5_nl;
  wire mux_2128_nl;
  wire mux_2130_nl;
  wire mux_2129_nl;
  wire mux_2131_nl;
  wire[39:0] attention_2_1_16_16_4_4_q_embed_mux1h_40_nl;
  wire attention_2_1_16_16_4_4_q_embed_or_nl;
  wire attention_2_1_16_16_4_4_q_embed_and_33_nl;
  wire not_4510_nl;
  wire mux_2156_nl;
  wire mux_2155_nl;
  wire nor_1240_nl;
  wire nor_1241_nl;
  wire nor_1242_nl;
  wire mux_2154_nl;
  wire nor_1243_nl;
  wire nor_1244_nl;
  wire[39:0] attention_2_1_16_16_4_4_q_embed_mux1h_41_nl;
  wire not_4483_nl;
  wire mux_2159_nl;
  wire mux_2158_nl;
  wire nor_1245_nl;
  wire[39:0] attention_2_1_16_16_4_4_q_embed_mux1h_42_nl;
  wire not_4482_nl;
  wire mux_2182_nl;
  wire mux_2181_nl;
  wire nor_1256_nl;
  wire[39:0] attention_2_1_16_16_4_4_q_embed_mux1h_43_nl;
  wire attention_2_1_16_16_4_4_q_embed_or_5_nl;
  wire attention_2_1_16_16_4_4_q_embed_and_35_nl;
  wire not_4511_nl;
  wire[39:0] attention_2_1_16_16_4_4_q_embed_mux1h_44_nl;
  wire not_4512_nl;
  wire mux_2198_nl;
  wire mux_2197_nl;
  wire nor_1272_nl;
  wire[39:0] attention_2_1_16_16_4_4_q_embed_mux1h_45_nl;
  wire not_4513_nl;
  wire mux_2204_nl;
  wire mux_2203_nl;
  wire nor_1283_nl;
  wire[39:0] attention_2_1_16_16_4_4_q_embed_mux1h_46_nl;
  wire not_4514_nl;
  wire mux_2210_nl;
  wire mux_2209_nl;
  wire nor_1294_nl;
  wire[39:0] attention_2_1_16_16_4_4_q_embed_mux1h_47_nl;
  wire attention_2_1_16_16_4_4_q_embed_or_6_nl;
  wire attention_2_1_16_16_4_4_q_embed_and_37_nl;
  wire not_4515_nl;
  wire[39:0] attention_2_1_16_16_4_4_q_embed_mux1h_48_nl;
  wire not_4516_nl;
  wire mux_2226_nl;
  wire mux_2225_nl;
  wire nor_1310_nl;
  wire[1:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_95_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_96_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_APPLY_ROTARY_POS_EMB_LOOP_6_or_7_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux_97_nl;
  wire[7:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_98_nl;
  wire[23:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_99_nl;
  wire[7:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_100_nl;
  wire[7:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux_101_nl;
  wire signed [55:0] nl_APPLY_ROTARY_POS_EMB_LOOP_6_mul_sgnd;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_and_35_nl;
  wire GEMM_3D_FLOAT_LOOP_3_not_28_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_and_34_nl;
  wire GEMM_3D_FLOAT_LOOP_3_not_27_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_and_33_nl;
  wire GEMM_3D_FLOAT_LOOP_3_not_26_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_and_32_nl;
  wire GEMM_3D_FLOAT_LOOP_3_not_25_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_and_31_nl;
  wire GEMM_3D_FLOAT_LOOP_3_not_24_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_and_30_nl;
  wire GEMM_3D_FLOAT_LOOP_3_not_23_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_and_29_nl;
  wire GEMM_3D_FLOAT_LOOP_3_not_22_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_and_28_nl;
  wire GEMM_3D_FLOAT_LOOP_3_not_21_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_and_27_nl;
  wire GEMM_3D_FLOAT_LOOP_3_not_20_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_and_26_nl;
  wire GEMM_3D_FLOAT_LOOP_3_not_19_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_and_25_nl;
  wire GEMM_3D_FLOAT_LOOP_3_not_18_nl;
  wire[39:0] GEMM_3D_FLOAT_LOOP_3_and_24_nl;
  wire GEMM_3D_FLOAT_LOOP_3_not_17_nl;
  wire mux_2237_nl;
  wire mux_1543_nl;
  wire mux_2248_nl;
  wire nor_1319_nl;
  wire mux_2250_nl;
  wire mux_2249_nl;
  wire mux_2258_nl;
  wire mux_2257_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_nl;
  wire not_4589_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_44_nl;
  wire not_4590_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_36_nl;
  wire not_4591_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_45_nl;
  wire not_4592_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_37_nl;
  wire not_4593_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_46_nl;
  wire not_4594_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_38_nl;
  wire not_4595_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_47_nl;
  wire not_4596_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_39_nl;
  wire not_4597_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_48_nl;
  wire not_4598_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_40_nl;
  wire not_4599_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_49_nl;
  wire not_4600_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_41_nl;
  wire not_4601_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_50_nl;
  wire not_4602_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_42_nl;
  wire not_4603_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_51_nl;
  wire not_4604_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_43_nl;
  wire not_4605_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_52_nl;
  wire not_4606_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_44_nl;
  wire not_4607_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_53_nl;
  wire not_4608_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_45_nl;
  wire not_4609_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_54_nl;
  wire not_4610_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_46_nl;
  wire not_4611_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_55_nl;
  wire not_4612_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_47_nl;
  wire not_4613_nl;
  wire[7:0] attention_2_1_16_16_4_4_k_proj_re_mux_56_nl;
  wire not_5055_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux_60_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux_61_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux_62_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux_63_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux_64_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux_65_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux_66_nl;
  wire attention_2_1_16_16_4_4_k_proj_re_mux_67_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_48_nl;
  wire not_4615_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_57_nl;
  wire not_4616_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_49_nl;
  wire not_4617_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_58_nl;
  wire not_4618_nl;
  wire[23:0] attention_2_1_16_16_4_4_v_proj_re_mux_50_nl;
  wire not_4619_nl;
  wire[15:0] attention_2_1_16_16_4_4_k_proj_re_mux_59_nl;
  wire not_4620_nl;
  wire output_and_35_nl;
  wire output_and_39_nl;
  wire output_and_43_nl;
  wire output_and_47_nl;
  wire output_and_51_nl;
  wire output_and_55_nl;
  wire output_and_59_nl;
  wire output_and_63_nl;
  wire output_and_61_nl;
  wire output_and_57_nl;
  wire output_and_53_nl;
  wire output_and_49_nl;
  wire output_and_45_nl;
  wire output_and_41_nl;
  wire output_and_37_nl;
  wire output_and_33_nl;
  wire or_1659_nl;
  wire nand_298_nl;
  wire or_1661_nl;
  wire nand_299_nl;
  wire or_1663_nl;
  wire nand_300_nl;
  wire or_1665_nl;
  wire nand_301_nl;
  wire or_1669_nl;
  wire or_1671_nl;
  wire[40:0] compute_sqrt_1_for_acc_1_nl;
  wire[41:0] nl_compute_sqrt_1_for_acc_1_nl;
  wire or_1860_nl;
  wire[40:0] compute_sqrt_for_acc_1_nl;
  wire[41:0] nl_compute_sqrt_for_acc_1_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_and_1_nl;
  wire[40:0] QUANTIZE_ACTIVATION_LOOP_2_acc_4_nl;
  wire[41:0] nl_QUANTIZE_ACTIVATION_LOOP_2_acc_4_nl;
  wire QUANTIZE_ACTIVATION_LOOP_2_attention_abs_2_nand_nl;
  wire[38:0] attention_abs_2_mux_3_nl;
  wire[25:0] QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_nl;
  wire[26:0] nl_QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_nl;
  wire[23:0] operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux_32_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_3_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_1_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_4_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_2_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_5_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_3_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_6_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_4_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_7_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_5_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_8_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_6_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_9_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_7_nl;
  wire[23:0] operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_17_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_5_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_1_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_6_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_2_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_7_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_3_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_8_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_4_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_9_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_5_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_10_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_6_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_11_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_7_nl;
  wire[23:0] operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_17_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_mux_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_3_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_mux_1_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_4_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_mux_2_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_5_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_mux_3_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_6_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_mux_4_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_7_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_mux_5_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_8_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_mux_6_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_9_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_mux_7_nl;
  wire[23:0] APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_1_nl;
  wire[7:0] APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_7_nl;
  wire[7:0] APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_25_nl;
  wire[23:0] APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_6_nl;
  wire[2:0] APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_26_nl;
  wire[2:0] APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_27_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_28_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_16_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_17_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_18_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_19_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_20_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_21_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_22_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_23_nl;
  wire nand_378_nl;
  wire[55:0] APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_nl;
  wire[56:0] nl_APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_nl;
  wire[55:0] APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_nl;
  wire[56:0] nl_APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_nl;
  wire or_3014_nl;
  wire or_3017_nl;
  wire or_3019_nl;
  wire or_3021_nl;
  wire or_3022_nl;
  wire or_3023_nl;
  wire or_3024_nl;
  wire or_3025_nl;
  wire or_3027_nl;
  wire or_3028_nl;
  wire or_3029_nl;
  wire or_3030_nl;
  wire SF_LOOP_3_and_nl;
  wire[23:0] operator_40_24_true_AC_TRN_AC_WRAP_acc_nl;
  wire[24:0] nl_operator_40_24_true_AC_TRN_AC_WRAP_acc_nl;
  wire[40:0] QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_nl;
  wire[41:0] nl_QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_nl;
  wire QUANTIZE_ACTIVATION_LOOP_2_1_attention_abs_6_nand_nl;
  wire[38:0] attention_abs_6_mux_3_nl;
  wire[25:0] QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_nl;
  wire[26:0] nl_QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_nl;
  wire[23:0] operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_mux_32_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_3_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_1_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_4_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_2_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_5_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_3_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_6_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_4_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_7_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_5_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_8_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_6_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_9_nl;
  wire LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_7_nl;
  wire[2:0] CACHE_UPDATE_LOOP_2_1_acc_2_nl;
  wire[3:0] nl_CACHE_UPDATE_LOOP_2_1_acc_2_nl;
  wire[40:0] attention_max_attn_fixed_t_1_acc_1_nl;
  wire[41:0] nl_attention_max_attn_fixed_t_1_acc_1_nl;
  wire[2:0] CACHE_UPDATE_LOOP_2_acc_2_nl;
  wire[3:0] nl_CACHE_UPDATE_LOOP_2_acc_2_nl;
  wire[40:0] SOFTMAX_LOOP_3_acc_3_nl;
  wire[41:0] nl_SOFTMAX_LOOP_3_acc_3_nl;
  wire mux_819_nl;
  wire mux_817_nl;
  wire mux_831_nl;
  wire mux_830_nl;
  wire mux_829_nl;
  wire mux_828_nl;
  wire mux_827_nl;
  wire nand_257_nl;
  wire or_1090_nl;
  wire mux_826_nl;
  wire mux_823_nl;
  wire mux_822_nl;
  wire mux_835_nl;
  wire mux_833_nl;
  wire mux_837_nl;
  wire and_1498_nl;
  wire nor_897_nl;
  wire and_337_nl;
  wire mux_858_nl;
  wire mux_867_nl;
  wire nand_262_nl;
  wire mux_866_nl;
  wire and_344_nl;
  wire or_3142_nl;
  wire mux_865_nl;
  wire or_1827_nl;
  wire mux_904_nl;
  wire nand_44_nl;
  wire mux_903_nl;
  wire mux_953_nl;
  wire or_3149_nl;
  wire or_3150_nl;
  wire nor_923_nl;
  wire nand_264_nl;
  wire or_1910_nl;
  wire or_1912_nl;
  wire or_3073_nl;
  wire mux_1026_nl;
  wire mux_1028_nl;
  wire or_1976_nl;
  wire or_1974_nl;
  wire mux_1149_nl;
  wire mux_1148_nl;
  wire mux_1162_nl;
  wire mux_1161_nl;
  wire mux_1160_nl;
  wire mux_1159_nl;
  wire mux_1158_nl;
  wire mux_1157_nl;
  wire mux_1156_nl;
  wire mux_1155_nl;
  wire mux_1154_nl;
  wire mux_1153_nl;
  wire mux_1152_nl;
  wire mux_1249_nl;
  wire mux_1311_nl;
  wire or_2235_nl;
  wire mux_1313_nl;
  wire nor_930_nl;
  wire mux_1312_nl;
  wire and_443_nl;
  wire mux_1400_nl;
  wire mux_1399_nl;
  wire mux_1398_nl;
  wire mux_1396_nl;
  wire and_1616_nl;
  wire mux_1395_nl;
  wire mux_1394_nl;
  wire or_2296_nl;
  wire mux_1406_nl;
  wire or_2309_nl;
  wire mux_1405_nl;
  wire mux_1404_nl;
  wire or_1049_nl;
  wire or_2322_nl;
  wire mux_1422_nl;
  wire and_1303_nl;
  wire mux_1425_nl;
  wire mux_1424_nl;
  wire mux_1423_nl;
  wire mux_1427_nl;
  wire or_2328_nl;
  wire mux_1436_nl;
  wire nor_938_nl;
  wire mux_1435_nl;
  wire nor_939_nl;
  wire mux_1450_nl;
  wire mux_1449_nl;
  wire mux_137_nl;
  wire mux_1942_nl;
  wire nor_946_nl;
  wire mux_1944_nl;
  wire or_2744_nl;
  wire mux_2035_nl;
  wire or_2746_nl;
  wire mux_2066_nl;
  wire mux_2085_nl;
  wire or_2784_nl;
  wire mux_2113_nl;
  wire mux_2112_nl;
  wire mux_2111_nl;
  wire nor_953_nl;
  wire nor_954_nl;
  wire nor_955_nl;
  wire mux_2110_nl;
  wire or_2833_nl;
  wire nor_956_nl;
  wire mux_2115_nl;
  wire mux_2117_nl;
  wire nor_957_nl;
  wire mux_2118_nl;
  wire mux_2152_nl;
  wire mux_2151_nl;
  wire mux_2150_nl;
  wire mux_2149_nl;
  wire mux_2148_nl;
  wire mux_2147_nl;
  wire nand_286_nl;
  wire or_2872_nl;
  wire mux_2145_nl;
  wire nand_101_nl;
  wire or_2869_nl;
  wire mux_2144_nl;
  wire or_2868_nl;
  wire mux_2143_nl;
  wire mux_2142_nl;
  wire or_2866_nl;
  wire mux_2175_nl;
  wire mux_2174_nl;
  wire mux_2173_nl;
  wire mux_2172_nl;
  wire mux_2171_nl;
  wire mux_2170_nl;
  wire or_2901_nl;
  wire mux_2169_nl;
  wire mux_2168_nl;
  wire and_1544_nl;
  wire mux_2165_nl;
  wire mux_2164_nl;
  wire mux_2162_nl;
  wire mux_2161_nl;
  wire mux_2160_nl;
  wire or_2897_nl;
  wire or_2894_nl;
  wire or_2890_nl;
  wire mux_2251_nl;
  wire and_1546_nl;
  wire nor_968_nl;
  wire or_3055_nl;
  wire or_3058_nl;
  wire mux_2255_nl;
  wire mux_2254_nl;
  wire mux_2253_nl;
  wire or_1418_nl;
  wire nand_295_nl;
  wire mux_2259_nl;
  wire and_1550_nl;
  wire nor_969_nl;
  wire mux_869_nl;
  wire mux_868_nl;
  wire mux_1010_nl;
  wire mux_1009_nl;
  wire mux_1008_nl;
  wire mux_1007_nl;
  wire nor_999_nl;
  wire mux_1006_nl;
  wire mux_1005_nl;
  wire nand_322_nl;
  wire nor_1001_nl;
  wire mux_1004_nl;
  wire mux_1003_nl;
  wire or_1952_nl;
  wire or_1950_nl;
  wire mux_1002_nl;
  wire mux_1001_nl;
  wire nand_323_nl;
  wire mux_999_nl;
  wire mux_998_nl;
  wire nand_325_nl;
  wire mux_997_nl;
  wire or_1944_nl;
  wire mux_996_nl;
  wire mux_995_nl;
  wire mux_994_nl;
  wire mux_993_nl;
  wire or_1943_nl;
  wire mux_992_nl;
  wire mux_991_nl;
  wire or_1940_nl;
  wire mux_990_nl;
  wire mux_989_nl;
  wire mux_988_nl;
  wire mux_987_nl;
  wire or_1939_nl;
  wire or_1938_nl;
  wire or_1937_nl;
  wire or_1934_nl;
  wire or_1933_nl;
  wire mux_986_nl;
  wire or_1932_nl;
  wire or_1931_nl;
  wire mux_1025_nl;
  wire mux_1024_nl;
  wire nor_1019_nl;
  wire mux_1023_nl;
  wire mux_1022_nl;
  wire mux_1021_nl;
  wire nor_1020_nl;
  wire nor_1021_nl;
  wire mux_1020_nl;
  wire nor_1022_nl;
  wire mux_1019_nl;
  wire nor_1023_nl;
  wire nor_1024_nl;
  wire mux_1032_nl;
  wire nand_49_nl;
  wire mux_1031_nl;
  wire mux_1030_nl;
  wire mux_1029_nl;
  wire mux_1078_nl;
  wire nor_1031_nl;
  wire nand_330_nl;
  wire mux_1076_nl;
  wire nor_1032_nl;
  wire nor_1033_nl;
  wire mux_1073_nl;
  wire or_2022_nl;
  wire mux_1077_nl;
  wire mux_1075_nl;
  wire or_2019_nl;
  wire mux_1088_nl;
  wire nand_52_nl;
  wire mux_1086_nl;
  wire mux_1085_nl;
  wire or_2038_nl;
  wire mux_1083_nl;
  wire mux_1082_nl;
  wire nand_332_nl;
  wire nand_51_nl;
  wire mux_1081_nl;
  wire nor_1035_nl;
  wire nor_1036_nl;
  wire or_2034_nl;
  wire mux_1080_nl;
  wire mux_1091_nl;
  wire or_2041_nl;
  wire mux_1090_nl;
  wire or_2039_nl;
  wire mux_1111_nl;
  wire or_2070_nl;
  wire mux_1110_nl;
  wire or_2068_nl;
  wire mux_1131_nl;
  wire mux_1130_nl;
  wire mux_1129_nl;
  wire mux_1128_nl;
  wire mux_1127_nl;
  wire mux_1126_nl;
  wire mux_1123_nl;
  wire mux_1121_nl;
  wire or_2095_nl;
  wire or_2110_nl;
  wire mux_1196_nl;
  wire mux_1195_nl;
  wire mux_1194_nl;
  wire mux_1193_nl;
  wire mux_1192_nl;
  wire mux_1191_nl;
  wire mux_1190_nl;
  wire mux_1189_nl;
  wire mux_1188_nl;
  wire mux_1186_nl;
  wire mux_1184_nl;
  wire mux_1182_nl;
  wire mux_1181_nl;
  wire mux_1180_nl;
  wire or_2121_nl;
  wire and_1593_nl;
  wire or_2132_nl;
  wire mux_1206_nl;
  wire mux_1205_nl;
  wire nor_1043_nl;
  wire and_1595_nl;
  wire mux_1204_nl;
  wire mux_1203_nl;
  wire or_2130_nl;
  wire mux_1202_nl;
  wire or_3166_nl;
  wire mux_1201_nl;
  wire or_2129_nl;
  wire mux_1200_nl;
  wire mux_1199_nl;
  wire or_2127_nl;
  wire mux_1198_nl;
  wire or_2126_nl;
  wire nor_1325_nl;
  wire mux_1273_nl;
  wire mux_1272_nl;
  wire mux_1271_nl;
  wire mux_1270_nl;
  wire or_2184_nl;
  wire nor_1050_nl;
  wire mux_1269_nl;
  wire mux_1268_nl;
  wire mux_1267_nl;
  wire mux_1266_nl;
  wire mux_1265_nl;
  wire nor_1326_nl;
  wire nor_1327_nl;
  wire mux_1264_nl;
  wire mux_1263_nl;
  wire nor_1328_nl;
  wire nor_1329_nl;
  wire mux_1262_nl;
  wire nor_1330_nl;
  wire nor_1331_nl;
  wire mux_1276_nl;
  wire mux_1275_nl;
  wire nor_1054_nl;
  wire nor_1055_nl;
  wire mux_1280_nl;
  wire or_3169_nl;
  wire mux_1279_nl;
  wire or_2199_nl;
  wire or_2198_nl;
  wire or_3170_nl;
  wire mux_1278_nl;
  wire or_2195_nl;
  wire mux_1277_nl;
  wire or_2193_nl;
  wire mux_1284_nl;
  wire mux_1283_nl;
  wire and_601_nl;
  wire nor_1060_nl;
  wire mux_1282_nl;
  wire or_2203_nl;
  wire nor_1102_nl;
  wire and_1635_nl;
  wire mux_1402_nl;
  wire mux_1401_nl;
  wire nor_1099_nl;
  wire nor_1100_nl;
  wire nor_1101_nl;
  wire mux_1409_nl;
  wire mux_1408_nl;
  wire mux_1407_nl;
  wire mux_1448_nl;
  wire and_1642_nl;
  wire mux_1447_nl;
  wire nor_1111_nl;
  wire mux_1446_nl;
  wire mux_1445_nl;
  wire mux_1444_nl;
  wire mux_1443_nl;
  wire mux_1442_nl;
  wire and_1644_nl;
  wire mux_1464_nl;
  wire nor_1118_nl;
  wire nor_1119_nl;
  wire mux_1463_nl;
  wire nor_1120_nl;
  wire mux_1462_nl;
  wire nor_1121_nl;
  wire mux_1461_nl;
  wire or_2363_nl;
  wire or_2362_nl;
  wire mux_1460_nl;
  wire mux_1459_nl;
  wire nor_1122_nl;
  wire nor_1123_nl;
  wire mux_1458_nl;
  wire nor_1124_nl;
  wire nor_1125_nl;
  wire mux_1474_nl;
  wire mux_1473_nl;
  wire nor_1129_nl;
  wire nor_1130_nl;
  wire and_1646_nl;
  wire mux_1472_nl;
  wire nor_1126_nl;
  wire mux_1471_nl;
  wire nor_1127_nl;
  wire nor_1128_nl;
  wire mux_1470_nl;
  wire mux_1469_nl;
  wire nor_1131_nl;
  wire nor_1132_nl;
  wire mux_1468_nl;
  wire mux_1467_nl;
  wire nor_1133_nl;
  wire nor_1134_nl;
  wire nor_1135_nl;
  wire mux_1586_nl;
  wire or_2499_nl;
  wire mux_1592_nl;
  wire nand_359_nl;
  wire mux_1594_nl;
  wire mux_2262_nl;
  wire mux_1595_nl;
  wire mux_1593_nl;
  wire mux_1596_nl;
  wire mux_1598_nl;
  wire mux_1597_nl;
  wire and_1659_nl;
  wire mux_1599_nl;
  wire mux_1607_nl;
  wire mux_1606_nl;
  wire nor_1160_nl;
  wire mux_1605_nl;
  wire nand_361_nl;
  wire nand_362_nl;
  wire mux_1604_nl;
  wire nor_1161_nl;
  wire mux_1603_nl;
  wire nor_1162_nl;
  wire nor_1163_nl;
  wire mux_1602_nl;
  wire nor_1164_nl;
  wire nor_1165_nl;
  wire mux_1601_nl;
  wire mux_1608_nl;
  wire and_1667_nl;
  wire mux_1610_nl;
  wire and_1666_nl;
  wire nor_1169_nl;
  wire and_1668_nl;
  wire mux_1609_nl;
  wire nor_1170_nl;
  wire nor_1171_nl;
  wire mux_1615_nl;
  wire mux_1614_nl;
  wire or_2541_nl;
  wire or_3189_nl;
  wire mux_2060_nl;
  wire or_2762_nl;
  wire mux_2069_nl;
  wire or_2768_nl;
  wire mux_2138_nl;
  wire and_1778_nl;
  wire mux_2137_nl;
  wire mux_2136_nl;
  wire or_1238_nl;
  wire nor_1234_nl;
  wire mux_2140_nl;
  wire mux_2135_nl;
  wire mux_2134_nl;
  wire mux_2133_nl;
  wire mux_2132_nl;
  wire and_1780_nl;
  wire nor_1261_nl;
  wire mux_2191_nl;
  wire mux_2186_nl;
  wire mux_2185_nl;
  wire mux_2184_nl;
  wire mux_2183_nl;
  wire nor_1299_nl;
  wire mux_2219_nl;
  wire mux_2214_nl;
  wire mux_2213_nl;
  wire mux_2212_nl;
  wire mux_2211_nl;
  wire GEMM_3D_FLOAT_LOOP_4_l_mux1h_6_nl;
  wire GEMM_3D_FLOAT_LOOP_4_l_mux1h_8_nl;
  wire QUANTIZE_ACTIVATION_LOOP_1_1_max_val_asn_GEMM_3D_FLOAT_LOOP_4_l_2_operator_40_24_true_AC_TRN_AC_WRAP_or_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_mux1h_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_or_nl;
  wire[3:0] compute_sqrt_for_acc_3_nl;
  wire[4:0] nl_compute_sqrt_for_acc_3_nl;
  wire RMS_NORM_LOOP_2_and_35_nl;
  wire nor_658_nl;
  wire RMS_NORM_LOOP_2_2_and_35_nl;
  wire mux_1260_nl;
  wire mux_1259_nl;
  wire mux_1258_nl;
  wire mux_1257_nl;
  wire mux_1256_nl;
  wire mux_1255_nl;
  wire mux_1254_nl;
  wire mux_1253_nl;
  wire mux_1252_nl;
  wire or_2167_nl;
  wire mux_1251_nl;
  wire mux_1247_nl;
  wire mux_1246_nl;
  wire mux_1244_nl;
  wire mux_1243_nl;
  wire or_3075_nl;
  wire mux_1242_nl;
  wire mux_1241_nl;
  wire nor_374_nl;
  wire mux_1239_nl;
  wire or_2162_nl;
  wire mux_1261_nl;
  wire nor_1048_nl;
  wire and_1603_nl;
  wire and_1256_nl;
  wire and_1257_nl;
  wire mux_2247_nl;
  wire mux_2246_nl;
  wire nor_1318_nl;
  wire[39:0] CACHE_UPDATE_LOOP_3_mux_3_nl;
  wire and_369_nl;
  wire[2:0] TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_nl;
  wire[3:0] nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_nl;
  wire[2:0] CACHE_UPDATE_LOOP_3_acc_nl;
  wire[3:0] nl_CACHE_UPDATE_LOOP_3_acc_nl;
  wire[23:0] CACHE_UPDATE_LOOP_3_1_CACHE_UPDATE_LOOP_3_1_mux_nl;
  wire[23:0] CACHE_UPDATE_LOOP_3_1_mux_2_nl;
  wire[15:0] CACHE_UPDATE_LOOP_3_1_CACHE_UPDATE_LOOP_3_1_mux_1_nl;
  wire[15:0] CACHE_UPDATE_LOOP_3_1_mux_3_nl;
  wire[2:0] GEMM_3D_FLOAT_LOOP_4_1_acc_13_nl;
  wire[3:0] nl_GEMM_3D_FLOAT_LOOP_4_1_acc_13_nl;
  wire[2:0] GEMM_3D_FLOAT_LOOP_4_acc_nl;
  wire[3:0] nl_GEMM_3D_FLOAT_LOOP_4_acc_nl;
  wire mux_2299_nl;
  wire nor_1345_nl;
  wire nor_1346_nl;
  wire mux_2288_nl;
  wire nor_1378_nl;
  wire nor_1379_nl;
  wire mux_2292_nl;
  wire or_3261_nl;
  wire mux_2291_nl;
  wire mux_2290_nl;
  wire or_3235_nl;
  wire mux_2267_nl;
  wire mux_2266_nl;
  wire nor_1348_nl;
  wire mux_2268_nl;
  wire nor_1350_nl;
  wire mux_2270_nl;
  wire nand_394_nl;
  wire mux_2287_nl;
  wire nor_1368_nl;
  wire mux_2286_nl;
  wire nand_398_nl;
  wire nor_1369_nl;
  wire CACHE_UPDATE_LOOP_3_mux1h_6_nl;
  wire CACHE_UPDATE_LOOP_3_mux1h_7_nl;
  wire GEMM_3D_FLOAT_LOOP_1_GEMM_3D_FLOAT_LOOP_1_mux_2_nl;
  wire GEMM_3D_FLOAT_LOOP_1_GEMM_3D_FLOAT_LOOP_1_mux_3_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_APPLY_ROTARY_POS_EMB_LOOP_6_or_8_nl;
  wire[12:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_36_nl;
  wire[23:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_37_nl;
  wire[7:0] APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_38_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_39_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_40_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_41_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_42_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_43_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_44_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_45_nl;
  wire APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_46_nl;
  wire RMS_NORM_LOOP_1_1_and_14_nl;
  wire RMS_NORM_LOOP_1_1_mux1h_134_nl;
  wire[2:0] RMS_NORM_LOOP_1_1_and_15_nl;
  wire[2:0] RMS_NORM_LOOP_1_1_mux1h_135_nl;
  wire RMS_NORM_LOOP_1_1_mux1h_136_nl;
  wire[5:0] RMS_NORM_LOOP_1_1_mux1h_137_nl;
  wire[4:0] RMS_NORM_LOOP_1_1_mux1h_138_nl;
  wire[7:0] RMS_NORM_LOOP_1_1_mux1h_139_nl;
  wire[7:0] RMS_NORM_LOOP_1_1_mux1h_140_nl;
  wire[7:0] RMS_NORM_LOOP_1_1_mux1h_141_nl;
  wire RMS_NORM_LOOP_1_1_and_16_nl;
  wire RMS_NORM_LOOP_1_1_mux1h_142_nl;
  wire[14:0] RMS_NORM_LOOP_1_1_and_17_nl;
  wire[14:0] RMS_NORM_LOOP_1_1_mux1h_143_nl;
  wire[6:0] RMS_NORM_LOOP_1_1_and_18_nl;
  wire[6:0] RMS_NORM_LOOP_1_1_mux1h_144_nl;
  wire not_5114_nl;
  wire RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_3_nl;
  wire RMS_NORM_LOOP_1_1_mux1h_145_nl;
  wire RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_4_nl;
  wire RMS_NORM_LOOP_1_1_mux1h_146_nl;
  wire[1:0] RMS_NORM_LOOP_1_1_and_19_nl;
  wire[1:0] RMS_NORM_LOOP_1_1_mux1h_147_nl;
  wire RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_5_nl;
  wire RMS_NORM_LOOP_1_1_mux1h_148_nl;
  wire[1:0] RMS_NORM_LOOP_1_1_mux1h_149_nl;
  wire RMS_NORM_LOOP_1_1_and_20_nl;
  wire RMS_NORM_LOOP_1_1_mux1h_150_nl;
  wire RMS_NORM_LOOP_1_1_or_13_nl;
  wire RMS_NORM_LOOP_1_1_mux1h_151_nl;
  wire[1:0] RMS_NORM_LOOP_1_1_mux1h_152_nl;
  wire RMS_NORM_LOOP_1_1_or_14_nl;
  wire RMS_NORM_LOOP_1_1_mux1h_153_nl;
  wire[4:0] RMS_NORM_LOOP_1_1_mux1h_154_nl;
  wire RMS_NORM_LOOP_1_1_or_15_nl;
  wire TRANSPOSE_LAST_TWO_DIMS_LOOP_3_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_mux_2_nl;
  wire TRANSPOSE_LAST_TWO_DIMS_LOOP_3_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_mux_3_nl;
  wire[3:0] RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_mux_1_nl;
  wire RMS_NORM_LOOP_2_2_or_1_nl;
  wire mux_2300_nl;
  wire mux_2301_nl;
  wire mux_2302_nl;
  wire nor_1397_nl;
  wire mux_2303_nl;
  wire nor_1398_nl;
  wire and_2128_nl;
  wire[71:0] mul_3_nl;
  wire signed [92:0] nl_mul_3_nl;
  wire[52:0] RMS_NORM_LOOP_2_2_mux_28_nl;
  wire and_2129_nl;
  wire[1:0] operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_21_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_22_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_23_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_22_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_23_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_24_nl;
  wire operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_25_nl;
  wire[2:0] RMS_NORM_LOOP_2_2_mux_29_nl;
  wire RMS_NORM_LOOP_2_2_mux_30_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [55:0] nl_SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a;
  assign nl_SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a = {SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_55
      , SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_54_16 , 16'b0000000000000000};
  wire [39:0] nl_SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b;
  assign nl_SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b = {SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_39
      , SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_38_0};
  wire [71:0] nl_LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a;
  assign nl_LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a
      = {LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_71_48
      , LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_47_40
      , LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_39
      , LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_38
      , LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_37
      , LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_36
      , LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_35
      , LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_34
      , LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_33
      , LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_32
      , 32'b00000000000000000000000000000000};
  wire [59:0] nl_LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b;
  assign nl_LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b
      = {LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_59_39
      , LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_38_0};
  wire [39:0] nl_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a;
  assign nl_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a = {1'b0, signext_39_33({reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd
      , 15'b000000000000000 , reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd_1
      , 16'b0000000000000000})};
  wire [39:0] nl_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b;
  assign nl_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b = {operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_39
      , operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_38_35 , operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_34
      , operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_33_0};
  wire[1:0] CACHE_UPDATE_LOOP_3_1_qif_acc_nl;
  wire[2:0] nl_CACHE_UPDATE_LOOP_3_1_qif_acc_nl;
  wire [4:0] nl_CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_rg_addr;
  assign nl_CACHE_UPDATE_LOOP_3_1_qif_acc_nl = conv_u2u_1_2(reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd)
      + ({reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign CACHE_UPDATE_LOOP_3_1_qif_acc_nl = nl_CACHE_UPDATE_LOOP_3_1_qif_acc_nl[1:0];
  assign nl_CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_rg_addr = {CACHE_UPDATE_LOOP_3_1_qif_acc_nl
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1};
  wire [5:0] nl_LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_rg_addr;
  assign nl_LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_rg_addr
      = {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2};
  wire [5:0] nl_LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_rg_addr;
  assign nl_LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_rg_addr
      = {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2};
  wire [9:0] nl_APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_rg_addr;
  assign nl_APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_rg_addr
      = {8'b00110000 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1};
  wire [9:0] nl_APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_rg_addr;
  assign nl_APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_rg_addr
      = {8'b00110000 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1};
  wire [5:0] nl_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_rg_addr;
  assign nl_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_rg_addr
      = {reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2};
  wire [5:0] nl_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_rg_addr;
  assign nl_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_rg_addr
      = {reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1
      , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1};
  wire[1:0] CACHE_UPDATE_LOOP_3_qif_acc_nl;
  wire[2:0] nl_CACHE_UPDATE_LOOP_3_qif_acc_nl;
  wire [4:0] nl_CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_rg_addr;
  assign nl_CACHE_UPDATE_LOOP_3_qif_acc_nl = conv_u2u_1_2(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[1])
      + ({reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign CACHE_UPDATE_LOOP_3_qif_acc_nl = nl_CACHE_UPDATE_LOOP_3_qif_acc_nl[1:0];
  assign nl_CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_rg_addr = {CACHE_UPDATE_LOOP_3_qif_acc_nl
      , (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]) , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1};
  wire [31:0] nl_dut_core_strm_out_rsci_inst_strm_out_rsci_idat;
  assign nl_dut_core_strm_out_rsci_inst_strm_out_rsci_idat = {strm_out_rsci_idat_31_18
      , strm_out_rsci_idat_17_10 , strm_out_rsci_idat_9 , strm_out_rsci_idat_8 ,
      strm_out_rsci_idat_7 , strm_out_rsci_idat_6 , strm_out_rsci_idat_5 , strm_out_rsci_idat_4
      , strm_out_rsci_idat_3 , strm_out_rsci_idat_2 , 2'b00};
  wire  nl_dut_core_core_fsm_inst_compute_sqrt_for_C_15_tr0;
  assign nl_dut_core_core_fsm_inst_compute_sqrt_for_C_15_tr0 = ~ reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  wire  nl_dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0 = (LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_2[2])
      & (z_out_5[2]) & (z_out_3[2]);
  wire  nl_dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0;
  assign nl_dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0 = (z_out_3[2])
      & (z_out_4[2]) & (z_out_5[2]);
  wire  nl_dut_core_core_fsm_inst_RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0 = (reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      | reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1) & (z_out_3[2]);
  wire  nl_dut_core_core_fsm_inst_APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0;
  assign nl_dut_core_core_fsm_inst_APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0 = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1];
  wire  nl_dut_core_core_fsm_inst_APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0 = z_out_4[2];
  wire  nl_dut_core_core_fsm_inst_CACHE_UPDATE_LOOP_3_C_1_tr0;
  assign nl_dut_core_core_fsm_inst_CACHE_UPDATE_LOOP_3_C_1_tr0 = reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1
      & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1]);
  wire  nl_dut_core_core_fsm_inst_CACHE_UPDATE_LOOP_2_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_CACHE_UPDATE_LOOP_2_C_0_tr0 = ~(CACHE_UPDATE_LOOP_2_acc_2_itm_2_1
      | CACHE_UPDATE_LOOP_2_1_acc_2_itm_2_1);
  wire  nl_dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0;
  assign nl_dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0 = TRANSPOSE_LAST_TWO_DIMS_LOOP_3_k_2_0_sva_1[2];
  wire  nl_dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0 = ~ CACHE_UPDATE_LOOP_2_1_acc_2_itm_2_1;
  wire  nl_dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0 = z_out_5[2];
  wire  nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_3_C_1_tr0;
  assign nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_3_C_1_tr0 = ~ CACHE_UPDATE_LOOP_2_1_acc_2_itm_2_1;
  wire  nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_1_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_1_C_0_tr0 = z_out_5[2];
  wire  nl_dut_core_core_fsm_inst_SF_LOOP_3_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_SF_LOOP_3_C_0_tr0 = ~ CACHE_UPDATE_LOOP_2_1_acc_2_itm_2_1;
  wire  nl_dut_core_core_fsm_inst_SF_LOOP_1_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_SF_LOOP_1_C_0_tr0 = z_out_5[2];
  wire  nl_dut_core_core_fsm_inst_CM_LOOP_1_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_CM_LOOP_1_C_0_tr0 = z_out_3[2];
  wire  nl_dut_core_core_fsm_inst_SOFTMAX_LOOP_3_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_SOFTMAX_LOOP_3_C_0_tr0 = ~ reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  wire  nl_dut_core_core_fsm_inst_SOFTMAX_LOOP_4_C_2_tr0;
  assign nl_dut_core_core_fsm_inst_SOFTMAX_LOOP_4_C_2_tr0 = ~ reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  wire  nl_dut_core_core_fsm_inst_SOFTMAX_LOOP_5_C_19_tr0;
  assign nl_dut_core_core_fsm_inst_SOFTMAX_LOOP_5_C_19_tr0 = ~ reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  wire  nl_dut_core_core_fsm_inst_SOFTMAX_LOOP_1_C_1_tr0;
  assign nl_dut_core_core_fsm_inst_SOFTMAX_LOOP_1_C_1_tr0 = z_out_5[2];
  wire  nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0;
  assign nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0 = ~ reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  wire  nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0;
  assign nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0 = z_out_4[2];
  wire  nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0 = z_out_5[2];
  wire  nl_dut_core_core_fsm_inst_ATTN_2D_LOOP_3_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_ATTN_2D_LOOP_3_C_0_tr0 = z_out_5[2];
  wire  nl_dut_core_core_fsm_inst_ATTN_2D_LOOP_2_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_ATTN_2D_LOOP_2_C_0_tr0 = z_out_4[2];
  wire  nl_dut_core_core_fsm_inst_compute_sqrt_1_for_C_15_tr0;
  assign nl_dut_core_core_fsm_inst_compute_sqrt_1_for_C_15_tr0 = ~ reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  wire  nl_dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0;
  assign nl_dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0 = z_out_5[2];
  wire  nl_dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0;
  assign nl_dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0 = z_out_4[2];
  mgc_div #(.width_a(32'sd56),
  .width_b(32'sd40),
  .signd(32'sd1)) SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp (
      .a(nl_SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a[55:0]),
      .b(nl_SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b[39:0]),
      .z(SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z)
    );
  mgc_div #(.width_a(32'sd72),
  .width_b(32'sd60),
  .signd(32'sd1)) LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp
      (
      .a(nl_LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a[71:0]),
      .b(nl_LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b[59:0]),
      .z(LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z)
    );
  mgc_div #(.width_a(32'sd40),
  .width_b(32'sd40),
  .signd(32'sd1)) operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp (
      .a(nl_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a[39:0]),
      .b(nl_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b[39:0]),
      .z(operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z)
    );
  dutmgc_rom_33_32_20_1  CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_rg
      (
      .addr(nl_CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_rg_addr[4:0]),
      .data_out(CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_sdt)
    );
  dutmgc_rom_34_64_8_1  LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_rg
      (
      .addr(nl_LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_rg_addr[5:0]),
      .data_out(LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_itm)
    );
  dutmgc_rom_35_64_8_1  LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_rg
      (
      .addr(nl_LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_rg_addr[5:0]),
      .data_out(LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_itm)
    );
  dutmgc_rom_36_960_15_1  APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_rg
      (
      .addr(nl_APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_rg_addr[9:0]),
      .data_out(APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_itm)
    );
  dutmgc_rom_37_960_13_1  APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_rg
      (
      .addr(nl_APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_rg_addr[9:0]),
      .data_out(APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm)
    );
  dutmgc_rom_38_64_8_1  LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_rg
      (
      .addr(nl_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_rg_addr[5:0]),
      .data_out(LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm)
    );
  dutmgc_rom_39_64_8_1  LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_rg
      (
      .addr(nl_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_rg_addr[5:0]),
      .data_out(LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm)
    );
  dutmgc_rom_40_32_19_1  CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_rg (
      .addr(nl_CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_rg_addr[4:0]),
      .data_out(CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_itm)
    );
  dut_core_strm_in_rsci dut_core_strm_in_rsci_inst (
      .strm_in_rsc_dat(strm_in_rsc_dat),
      .strm_in_rsc_vld(strm_in_rsc_vld),
      .strm_in_rsc_rdy(strm_in_rsc_rdy),
      .strm_in_rsci_oswt(reg_strm_in_rsci_iswt0_cse),
      .strm_in_rsci_wen_comp(strm_in_rsci_wen_comp),
      .strm_in_rsci_idat_mxwt(strm_in_rsci_idat_mxwt)
    );
  dut_core_strm_out_rsci dut_core_strm_out_rsci_inst (
      .strm_out_rsc_dat(strm_out_rsc_dat),
      .strm_out_rsc_vld(strm_out_rsc_vld),
      .strm_out_rsc_rdy(strm_out_rsc_rdy),
      .strm_out_rsci_oswt(reg_strm_out_rsci_iswt0_cse),
      .strm_out_rsci_wen_comp(strm_out_rsci_wen_comp),
      .strm_out_rsci_idat(nl_dut_core_strm_out_rsci_inst_strm_out_rsci_idat[31:0])
    );
  dut_core_staller dut_core_staller_inst (
      .en(en),
      .core_wen1(core_wen1),
      .strm_in_rsci_wen_comp(strm_in_rsci_wen_comp),
      .strm_out_rsci_wen_comp(strm_out_rsci_wen_comp),
      .attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1(attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1)
    );
  dut_core_wait_dp dut_core_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .rms_norm_16_div_cmp_z(rms_norm_16_div_cmp_z),
      .core_wen1(core_wen1),
      .rms_norm_16_div_cmp_z_oreg(rms_norm_16_div_cmp_z_oreg)
    );
  dut_core_core_fsm dut_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1(attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1),
      .fsm_output(fsm_output),
      .for_for_C_2_tr0(for_for_and_tmp),
      .compute_sqrt_for_C_15_tr0(nl_dut_core_core_fsm_inst_compute_sqrt_for_C_15_tr0),
      .RMS_NORM_LOOP_2_C_4_tr0(and_37_cse),
      .QUANTIZE_ACTIVATION_LOOP_3_C_2_tr0(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4),
      .LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0(nl_dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_4_C_0_tr0),
      .LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0(nl_dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_3_C_1_tr0),
      .LINEAR_FORWARD_NO_MUL_LOOP_2_C_63_tr0(reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1),
      .RESHAPE_2D_TO_3D_LOOP_3_C_0_tr0(CACHE_UPDATE_LOOP_1_and_tmp),
      .RESHAPE_2D_TO_3D_LOOP_2_C_0_tr0(RESHAPE_2D_TO_3D_LOOP_2_2_and_cse),
      .RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0(nl_dut_core_core_fsm_inst_RESHAPE_2D_TO_3D_LOOP_3_2_C_0_tr0),
      .RESHAPE_2D_TO_3D_LOOP_2_2_C_0_tr0(RESHAPE_2D_TO_3D_LOOP_2_2_and_cse),
      .APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0(nl_dut_core_core_fsm_inst_APPLY_ROTARY_POS_EMB_LOOP_6_C_2_tr0),
      .APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0(nl_dut_core_core_fsm_inst_APPLY_ROTARY_POS_EMB_LOOP_4_C_0_tr0),
      .CACHE_UPDATE_LOOP_3_C_1_tr0(nl_dut_core_core_fsm_inst_CACHE_UPDATE_LOOP_3_C_1_tr0),
      .CACHE_UPDATE_LOOP_2_C_0_tr0(nl_dut_core_core_fsm_inst_CACHE_UPDATE_LOOP_2_C_0_tr0),
      .CACHE_UPDATE_LOOP_1_C_0_tr0(CACHE_UPDATE_LOOP_1_and_tmp),
      .TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0(nl_dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_C_2_tr0),
      .TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0(nl_dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_2_C_0_tr0),
      .TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0(nl_dut_core_core_fsm_inst_TRANSPOSE_LAST_TWO_DIMS_LOOP_1_C_0_tr0),
      .GEMM_3D_FLOAT_LOOP_4_C_3_tr0(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1),
      .GEMM_3D_FLOAT_LOOP_3_C_1_tr0(nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_3_C_1_tr0),
      .GEMM_3D_FLOAT_LOOP_1_C_0_tr0(nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_1_C_0_tr0),
      .SF_LOOP_3_C_0_tr0(nl_dut_core_core_fsm_inst_SF_LOOP_3_C_0_tr0),
      .SF_LOOP_1_C_0_tr0(nl_dut_core_core_fsm_inst_SF_LOOP_1_C_0_tr0),
      .CM_LOOP_1_C_0_tr0(nl_dut_core_core_fsm_inst_CM_LOOP_1_C_0_tr0),
      .SOFTMAX_LOOP_3_C_0_tr0(nl_dut_core_core_fsm_inst_SOFTMAX_LOOP_3_C_0_tr0),
      .SOFTMAX_LOOP_4_C_2_tr0(nl_dut_core_core_fsm_inst_SOFTMAX_LOOP_4_C_2_tr0),
      .SOFTMAX_LOOP_5_C_19_tr0(nl_dut_core_core_fsm_inst_SOFTMAX_LOOP_5_C_19_tr0),
      .SOFTMAX_LOOP_1_C_1_tr0(nl_dut_core_core_fsm_inst_SOFTMAX_LOOP_1_C_1_tr0),
      .GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0(nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_4_1_C_3_tr0),
      .GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0(nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_3_1_C_1_tr0),
      .GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0(nl_dut_core_core_fsm_inst_GEMM_3D_FLOAT_LOOP_1_1_C_0_tr0),
      .ATTN_2D_LOOP_3_C_0_tr0(nl_dut_core_core_fsm_inst_ATTN_2D_LOOP_3_C_0_tr0),
      .ATTN_2D_LOOP_2_C_0_tr0(nl_dut_core_core_fsm_inst_ATTN_2D_LOOP_2_C_0_tr0),
      .RMS_NORM_LOOP_1_2_C_2_tr0(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4),
      .compute_sqrt_1_for_C_15_tr0(nl_dut_core_core_fsm_inst_compute_sqrt_1_for_C_15_tr0),
      .RMS_NORM_LOOP_2_2_C_4_tr0(and_37_cse),
      .QUANTIZE_ACTIVATION_LOOP_3_1_C_2_tr0(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4),
      .LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0(nl_dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_4_3_C_0_tr0),
      .LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0(nl_dut_core_core_fsm_inst_LINEAR_FORWARD_NO_MUL_LOOP_3_3_C_1_tr0),
      .LINEAR_FORWARD_NO_MUL_LOOP_2_3_C_31_tr0(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4),
      .for_1_for_C_1_tr0(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4)
    );
  assign attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1;
  assign for_1_for_and_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 &
      (~(or_dcpl_961 | (~((fsm_output[5]) & (fsm_output[3]))) | or_1984_cse));
  assign attention_2_1_16_16_4_4_attn_output_and_4_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & and_dcpl_187;
  assign nand_302_cse = ~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva);
  assign nand_303_tmp = ~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva);
  assign attention_2_1_16_16_4_4_attn_output_and_14_cse = nand_303_tmp & and_dcpl_187;
  assign attention_2_1_16_16_4_4_attn_output_and_13_cse = (~ nand_303_tmp) & and_dcpl_187;
  assign nand_304_tmp = ~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva);
  assign attention_2_1_16_16_4_4_attn_output_and_16_cse = nand_304_tmp & and_dcpl_187;
  assign attention_2_1_16_16_4_4_attn_output_and_15_cse = (~ nand_304_tmp) & and_dcpl_187;
  assign nand_305_tmp = ~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva);
  assign attention_2_1_16_16_4_4_attn_output_and_18_cse = nand_305_tmp & and_dcpl_187;
  assign attention_2_1_16_16_4_4_attn_output_and_17_cse = (~ nand_305_tmp) & and_dcpl_187;
  assign and_1481_nl = (((fsm_output[2]) & (fsm_output[6])) | (fsm_output[7])) &
      (fsm_output[8]);
  assign mux_775_nl = MUX_s_1_2_2(and_1481_nl, mux_tmp_363, fsm_output[5]);
  assign or_1677_nl = (z_out_5[2]) | (~ (fsm_output[5])) | (fsm_output[2]);
  assign mux_774_nl = MUX_s_1_2_2(mux_tmp_363, nor_tmp_117, or_1677_nl);
  assign mux_776_nl = MUX_s_1_2_2(mux_775_nl, mux_774_nl, fsm_output[3]);
  assign or_1676_nl = (fsm_output[3]) | (~ (fsm_output[5])) | (fsm_output[2]);
  assign mux_773_nl = MUX_s_1_2_2(mux_tmp_363, nor_tmp_117, or_1676_nl);
  assign mux_777_nl = MUX_s_1_2_2(mux_776_nl, mux_773_nl, or_1732_cse);
  assign mux_778_nl = MUX_s_1_2_2(mux_777_nl, nor_tmp_117, fsm_output[4]);
  assign attention_2_1_16_16_4_4_attn_weights_and_36_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & mux_778_nl;
  assign attention_2_1_16_16_4_4_q_embed_and_5_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & and_dcpl_204;
  assign attention_2_1_16_16_4_4_q_embed_and_23_cse = (~ or_dcpl_991) & and_dcpl_204;
  assign attention_2_1_16_16_4_4_q_embed_and_24_cse = or_dcpl_991 & and_dcpl_204;
  assign attention_2_1_16_16_4_4_q_embed_mux_7_cse = MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_q_embed_2_0_3_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1, attention_2_1_16_16_4_4_q_embed_2_0_3_lpi_3,
      {(~ and_dcpl_204) , attention_2_1_16_16_4_4_q_embed_and_23_cse , attention_2_1_16_16_4_4_q_embed_and_24_cse});
  assign attention_2_1_16_16_4_4_q_embed_and_25_cse = (~ or_dcpl_995) & and_dcpl_204;
  assign attention_2_1_16_16_4_4_q_embed_and_26_cse = or_dcpl_995 & and_dcpl_204;
  assign attention_2_1_16_16_4_4_q_embed_mux_9_cse = MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_q_embed_3_0_0_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1, attention_2_1_16_16_4_4_q_embed_3_0_0_lpi_3,
      {(~ and_dcpl_204) , attention_2_1_16_16_4_4_q_embed_and_25_cse , attention_2_1_16_16_4_4_q_embed_and_26_cse});
  assign attention_2_1_16_16_4_4_q_embed_and_27_cse = (~ or_dcpl_997) & and_dcpl_204;
  assign attention_2_1_16_16_4_4_q_embed_and_28_cse = or_dcpl_997 & and_dcpl_204;
  assign attention_2_1_16_16_4_4_q_embed_mux_11_cse = MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_q_embed_3_0_1_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1, attention_2_1_16_16_4_4_q_embed_3_0_1_lpi_3,
      {(~ and_dcpl_204) , attention_2_1_16_16_4_4_q_embed_and_27_cse , attention_2_1_16_16_4_4_q_embed_and_28_cse});
  assign attention_2_1_16_16_4_4_q_embed_and_29_cse = (~ or_dcpl_999) & and_dcpl_204;
  assign attention_2_1_16_16_4_4_q_embed_and_30_cse = or_dcpl_999 & and_dcpl_204;
  assign attention_2_1_16_16_4_4_q_embed_mux_13_cse = MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_q_embed_3_0_2_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1, attention_2_1_16_16_4_4_q_embed_3_0_2_lpi_3,
      {(~ and_dcpl_204) , attention_2_1_16_16_4_4_q_embed_and_29_cse , attention_2_1_16_16_4_4_q_embed_and_30_cse});
  assign attention_2_1_16_16_4_4_q_embed_and_31_nl = (~ or_dcpl_1000) & and_dcpl_204;
  assign attention_2_1_16_16_4_4_q_embed_and_32_nl = or_dcpl_1000 & and_dcpl_204;
  assign attention_2_1_16_16_4_4_q_embed_mux_14_cse = MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_q_embed_3_0_3_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1, attention_2_1_16_16_4_4_q_embed_3_0_3_lpi_3,
      {(~ and_dcpl_204) , attention_2_1_16_16_4_4_q_embed_and_31_nl , attention_2_1_16_16_4_4_q_embed_and_32_nl});
  assign attention_2_1_16_16_4_4_v_proj_and_2_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & and_dcpl_207;
  assign nor_728_nl = ~((fsm_output[4]) | (fsm_output[7]));
  assign mux_781_nl = MUX_s_1_2_2(nor_728_nl, (fsm_output[7]), fsm_output[6]);
  assign mux_782_nl = MUX_s_1_2_2(mux_781_nl, and_dcpl_148, fsm_output[2]);
  assign mux_783_nl = MUX_s_1_2_2(mux_782_nl, nor_tmp_261, fsm_output[1]);
  assign and_1383_nl = (fsm_output[4]) & (fsm_output[7]);
  assign mux_779_nl = MUX_s_1_2_2(and_dcpl_148, and_1383_nl, fsm_output[2]);
  assign mux_780_nl = MUX_s_1_2_2(nor_tmp_261, mux_779_nl, fsm_output[1]);
  assign mux_784_nl = MUX_s_1_2_2(mux_783_nl, mux_780_nl, fsm_output[0]);
  assign and_1485_nl = or_1879_cse & (fsm_output[7]);
  assign mux_785_nl = MUX_s_1_2_2(mux_784_nl, and_1485_nl, fsm_output[3]);
  assign mux_786_nl = MUX_s_1_2_2(mux_785_nl, (fsm_output[7]), fsm_output[5]);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_and_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (mux_786_nl | (fsm_output[8]));
  assign apply_rotary_pos_emb_1_4_4_rotated_q_or_11_cse = (and_dcpl_186 & and_dcpl_209)
      | ((~ RESHAPE_2D_TO_3D_LOOP_2_2_and_cse) & and_dcpl_213);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_or_12_cse = (RESHAPE_2D_TO_3D_LOOP_2_2_and_cse
      & and_dcpl_213) | and_dcpl_216;
  assign or_1732_cse = (fsm_output[1:0]!=2'b00);
  assign mux_792_cse = MUX_s_1_2_2((fsm_output[7]), (~ (fsm_output[7])), fsm_output[6]);
  assign attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1 = MUX_v_24_16_2(attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_3_39_16, apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_39_16,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16, attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_3_39_16, attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_3_39_16, attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_3_39_16, attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_3_39_16, attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_3_39_16, attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_3_39_16, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign attention_2_1_16_16_4_4_q_proj_and_23_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & and_dcpl_240;
  assign RESHAPE_2D_TO_3D_LOOP_3_1_mux_13_cse = MUX_v_8_2_2((z_out_1[15:8]), LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8,
      or_dcpl_1011);
  assign RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_7 = MUX_s_1_2_2((z_out_1[7]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd,
      or_dcpl_1011);
  assign RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_6 = MUX_s_1_2_2((z_out_1[6]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1,
      or_dcpl_1011);
  assign RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_5 = MUX_s_1_2_2((z_out_1[5]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2,
      or_dcpl_1011);
  assign RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_4 = MUX_s_1_2_2((z_out_1[4]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3,
      or_dcpl_1011);
  assign RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_3 = MUX_s_1_2_2((z_out_1[3]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4,
      or_dcpl_1011);
  assign RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_2 = MUX_s_1_2_2((z_out_1[2]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5,
      or_dcpl_1011);
  assign RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_1 = MUX_s_1_2_2((z_out_1[1]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6,
      or_dcpl_1011);
  assign RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_0 = MUX_s_1_2_2((z_out_1[0]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7,
      or_dcpl_1011);
  assign and_274_nl = or_1732_cse & mux_tmp_121;
  assign mux_801_nl = MUX_s_1_2_2(and_274_nl, nor_tmp_28, or_2699_cse);
  assign nor_271_nl = ~(and_37_cse | (fsm_output[1:0]!=2'b01));
  assign mux_799_nl = MUX_s_1_2_2(nor_tmp_28, mux_tmp_121, nor_271_nl);
  assign mux_800_nl = MUX_s_1_2_2(nor_tmp_28, mux_799_nl, and_1762_cse);
  assign mux_802_nl = MUX_s_1_2_2(mux_801_nl, mux_800_nl, fsm_output[3]);
  assign mux_803_nl = MUX_s_1_2_2(mux_802_nl, nor_tmp_28, fsm_output[2]);
  assign mux_804_nl = MUX_s_1_2_2(mux_803_nl, (fsm_output[8]), fsm_output[7]);
  assign input_and_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & mux_804_nl;
  assign and_1555_cse = (fsm_output[0]) & (fsm_output[2]);
  assign or_1769_cse = (~ (fsm_output[5])) | (fsm_output[8]);
  assign or_1770_cse = (fsm_output[5]) | (~ (fsm_output[8]));
  assign and_1559_cse = (fsm_output[2:1]==2'b11);
  assign mux_806_cse = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[6]);
  assign nor_973_cse = ~((fsm_output[7:6]!=2'b00));
  assign or_270_cse = (~ (fsm_output[2])) | (fsm_output[4]);
  assign or_1767_cse = (~ (fsm_output[7])) | (fsm_output[5]) | (fsm_output[8]);
  assign or_1772_cse = (fsm_output[4]) | (fsm_output[7]) | (fsm_output[5]) | (fsm_output[8]);
  assign or_1775_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[5]) | (fsm_output[8]);
  assign or_1774_nl = (fsm_output[1]) | and_1555_cse | (fsm_output[7]) | (fsm_output[5])
      | (fsm_output[8]);
  assign mux_814_nl = MUX_s_1_2_2(or_1775_nl, or_1774_nl, fsm_output[4]);
  assign mux_815_nl = MUX_s_1_2_2(mux_814_nl, or_1772_cse, fsm_output[3]);
  assign mux_811_nl = MUX_s_1_2_2(or_1770_cse, or_1769_cse, fsm_output[7]);
  assign or_1771_nl = (fsm_output[2:0]!=3'b000) | mux_811_nl;
  assign mux_812_nl = MUX_s_1_2_2(or_1771_nl, or_1767_cse, fsm_output[4]);
  assign nand_41_nl = ~((fsm_output[4]) & (~(and_1559_cse | (~ (fsm_output[7])) |
      (fsm_output[5]) | (fsm_output[8]))));
  assign mux_813_nl = MUX_s_1_2_2(mux_812_nl, nand_41_nl, fsm_output[3]);
  assign mux_816_ssc = MUX_s_1_2_2(mux_815_nl, mux_813_nl, fsm_output[6]);
  assign and_303_ssc = (~ mux_tmp_836) & and_dcpl_270;
  assign compute_sqrt_guess_or_1_ssc = ((~ and_dcpl_290) & and_dcpl_272 & nor_777_cse
      & and_dcpl_209) | ((~ and_dcpl_292) & and_dcpl_226 & (~ (fsm_output[1])) &
      ((fsm_output[4]) ^ (fsm_output[5])) & (~((fsm_output[0]) | (fsm_output[3])))
      & and_dcpl_148);
  assign mux_838_nl = MUX_s_1_2_2(or_3185_cse, (~ and_1559_cse), fsm_output[3]);
  assign and_315_ssc = mux_838_nl & (~ (fsm_output[8])) & and_dcpl_279 & and_dcpl_148;
  assign or_1803_nl = (fsm_output[1]) | (~ (fsm_output[4])) | (fsm_output[7]) | (fsm_output[5])
      | (fsm_output[8]);
  assign mux_848_nl = MUX_s_1_2_2(or_1772_cse, mux_tmp_841, fsm_output[1]);
  assign mux_849_nl = MUX_s_1_2_2(or_1803_nl, mux_848_nl, fsm_output[3]);
  assign mux_845_nl = MUX_s_1_2_2((fsm_output[5]), or_1769_cse, fsm_output[7]);
  assign or_1802_nl = (fsm_output[4]) | mux_845_nl;
  assign mux_846_nl = MUX_s_1_2_2(or_1802_nl, mux_tmp_839, or_1732_cse);
  assign or_1799_nl = (~ (fsm_output[4])) | (~ (fsm_output[7])) | (fsm_output[5])
      | (fsm_output[8]);
  assign mux_847_nl = MUX_s_1_2_2(mux_846_nl, or_1799_nl, fsm_output[3]);
  assign mux_850_nl = MUX_s_1_2_2(mux_849_nl, mux_847_nl, fsm_output[6]);
  assign or_1798_nl = (~ (fsm_output[4])) | (fsm_output[7]) | (fsm_output[5]) | (fsm_output[8]);
  assign mux_842_nl = MUX_s_1_2_2(or_1798_nl, or_1772_cse, or_1732_cse);
  assign mux_843_nl = MUX_s_1_2_2(mux_842_nl, mux_tmp_841, fsm_output[3]);
  assign or_1792_nl = (fsm_output[1]) | (~ (fsm_output[4])) | (~ (fsm_output[7]))
      | (fsm_output[5]) | (fsm_output[8]);
  assign mux_840_nl = MUX_s_1_2_2(mux_tmp_839, or_1792_nl, fsm_output[3]);
  assign mux_844_nl = MUX_s_1_2_2(mux_843_nl, mux_840_nl, fsm_output[6]);
  assign mux_851_ssc = MUX_s_1_2_2(mux_850_nl, mux_844_nl, fsm_output[2]);
  assign nor_977_nl = ~((fsm_output[6]) | mux_tmp_836);
  assign and_1561_nl = (~((fsm_output[2:1]==2'b11))) & (fsm_output[4]);
  assign mux_852_nl = MUX_s_1_2_2(nor_tmp_285, and_1561_nl, fsm_output[3]);
  assign and_1562_nl = (fsm_output[6]) & mux_852_nl;
  assign mux_853_nl = MUX_s_1_2_2(nor_977_nl, and_1562_nl, fsm_output[7]);
  assign and_321_ssc = mux_853_nl & and_dcpl_1;
  assign and_1474_cse = (fsm_output[1:0]==2'b11);
  assign mux_854_nl = MUX_s_1_2_2(and_1762_cse, (~ or_tmp_755), fsm_output[6]);
  assign and_329_ssc = mux_854_nl & and_dcpl_295;
  assign and_334_ssc = (~((~(nand_197_cse & (fsm_output[3:2]==2'b00))) & (fsm_output[4])))
      & and_dcpl_298;
  assign and_336_ssc = and_dcpl_206 & and_dcpl_302;
  assign or_1812_nl = (fsm_output[5]) | (fsm_output[4]) | (~ (fsm_output[8]));
  assign mux_855_nl = MUX_s_1_2_2(or_1770_cse, or_1812_nl, fsm_output[3]);
  assign nor_979_nl = ~((fsm_output[6]) | mux_855_nl);
  assign and_1564_nl = (fsm_output[6]) & (fsm_output[3]) & (fsm_output[5]) & (~ or_tmp_757);
  assign mux_856_ssc = MUX_s_1_2_2(nor_979_nl, and_1564_nl, fsm_output[7]);
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_2_or_1_cse = and_dcpl_257 | and_dcpl_265;
  assign mux_859_nl = MUX_s_1_2_2(mux_tmp_87, and_1771_cse, fsm_output[1]);
  assign mux_860_nl = MUX_s_1_2_2(mux_859_nl, nor_tmp_289, fsm_output[0]);
  assign mux_861_nl = MUX_s_1_2_2(mux_860_nl, (fsm_output[4]), fsm_output[3]);
  assign and_339_ssc = (~ mux_861_nl) & and_dcpl_298;
  assign mux_863_nl = MUX_s_1_2_2((~ nor_tmp_291), nor_tmp_282, fsm_output[5]);
  assign mux_864_nl = MUX_s_1_2_2(mux_863_nl, mux_tmp_91, fsm_output[3]);
  assign and_343_itm = (~ mux_864_nl) & and_dcpl_308;
  assign rms_norm_16_div_cmp_b = {reg_rms_norm_16_div_cmp_b_ftd_59_38 , reg_rms_norm_16_div_cmp_b_ftd_37_0
      , reg_rms_norm_16_div_cmp_b_ftd_1};
  assign rms_norm_16_div_cmp_a = {reg_rms_norm_16_div_cmp_a_ftd , reg_rms_norm_16_div_cmp_a_ftd_1_15_8
      , reg_rms_norm_16_div_cmp_a_ftd_1_7 , reg_rms_norm_16_div_cmp_a_ftd_1_6 , reg_rms_norm_16_div_cmp_a_ftd_1_5
      , reg_rms_norm_16_div_cmp_a_ftd_1_4 , reg_rms_norm_16_div_cmp_a_ftd_1_3 , reg_rms_norm_16_div_cmp_a_ftd_1_2
      , reg_rms_norm_16_div_cmp_a_ftd_1_1 , reg_rms_norm_16_div_cmp_a_ftd_1_0 , 32'b00000000000000000000000000000000};
  assign and_362_ssc = and_dcpl_322 & and_dcpl_319 & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      & (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign nor_907_nl = ~((fsm_output[3]) | (fsm_output[5]) | (fsm_output[0]) | (fsm_output[1])
      | (fsm_output[2]) | (fsm_output[4]) | (~ (fsm_output[8])));
  assign mux_873_nl = MUX_s_1_2_2((fsm_output[8]), nor_907_nl, fsm_output[6]);
  assign mux_870_nl = MUX_s_1_2_2(or_tmp_757, (fsm_output[8]), fsm_output[5]);
  assign or_85_nl = nor_646_cse | (fsm_output[8]);
  assign mux_871_nl = MUX_s_1_2_2(mux_870_nl, or_85_nl, fsm_output[3]);
  assign mux_872_nl = MUX_s_1_2_2(mux_871_nl, (fsm_output[8]), fsm_output[6]);
  assign mux_874_nl = MUX_s_1_2_2((~ mux_873_nl), mux_872_nl, fsm_output[7]);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_and_3_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & mux_874_nl;
  assign nor_294_nl = ~((~ (fsm_output[4])) | reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      | reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      | (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1));
  assign mux_876_nl = MUX_s_1_2_2(nor_tmp_117, mux_tmp_363, nor_294_nl);
  assign mux_877_nl = MUX_s_1_2_2(and_1455_cse, mux_876_nl, fsm_output[0]);
  assign mux_878_nl = MUX_s_1_2_2(mux_877_nl, nor_tmp_117, or_1835_cse);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_and_6_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & mux_878_nl;
  assign or_1840_nl = (~ (fsm_output[4])) | reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      | reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 | (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd)
      | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign mux_880_nl = MUX_s_1_2_2(mux_tmp_363, nor_tmp_117, or_1840_nl);
  assign mux_881_nl = MUX_s_1_2_2(and_1455_cse, mux_880_nl, fsm_output[0]);
  assign mux_882_nl = MUX_s_1_2_2(mux_881_nl, nor_tmp_117, or_1835_cse);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_and_7_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & mux_882_nl;
  assign nor_301_nl = ~((~ (fsm_output[4])) | reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      | reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 | (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd)
      | (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1));
  assign mux_884_nl = MUX_s_1_2_2(nor_tmp_117, mux_tmp_363, nor_301_nl);
  assign mux_885_nl = MUX_s_1_2_2(and_1455_cse, mux_884_nl, fsm_output[0]);
  assign mux_886_nl = MUX_s_1_2_2(mux_885_nl, nor_tmp_117, or_1835_cse);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_and_8_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & mux_886_nl;
  assign or_1848_cse = (~ (fsm_output[1])) | (~ (fsm_output[0])) | (fsm_output[8]);
  assign or_1851_cse = (fsm_output[5]) | (fsm_output[8]);
  assign nor_305_cse = ~((fsm_output[5]) | (~ (fsm_output[1])) | (~ (fsm_output[0])));
  assign ATTN_2D_LOOP_3_mux_16_itm = MUX_s_1_16_2((apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2[39]),
      (attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2[39]), (attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2[39]),
      attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_39, (attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2[39]),
      (attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2[39]), (attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2[39]),
      (attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2[39]), (attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2[39]),
      (attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2[39]), (attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2[39]),
      (attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2[39]), (attention_2_1_16_16_4_4_attn_output_3_0_0_sva_2[39]),
      (attention_2_1_16_16_4_4_attn_output_3_0_1_sva_2[39]), (attention_2_1_16_16_4_4_attn_output_3_0_2_sva_2[39]),
      (attention_2_1_16_16_4_4_attn_output_3_0_3_sva_2[39]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign ATTN_2D_LOOP_3_mux_17_itm = MUX_v_39_16_2((apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2[38:0]),
      (attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2[38:0]), (attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2[38:0]),
      attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_38_0, (attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2[38:0]),
      (attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2[38:0]), (attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2[38:0]),
      (attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2[38:0]), (attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2[38:0]),
      (attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2[38:0]), (attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2[38:0]),
      (attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2[38:0]), (attention_2_1_16_16_4_4_attn_output_3_0_0_sva_2[38:0]),
      (attention_2_1_16_16_4_4_attn_output_3_0_1_sva_2[38:0]), (attention_2_1_16_16_4_4_attn_output_3_0_2_sva_2[38:0]),
      (attention_2_1_16_16_4_4_attn_output_3_0_3_sva_2[38:0]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign or_1880_cse = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 | reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign and_28_cse = (input_0_0_sva_2[39]) & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign or_1879_cse = (fsm_output[4]) | (fsm_output[6]);
  assign or_1867_cse = (~ (fsm_output[1])) | (fsm_output[4]);
  assign GEMM_3D_FLOAT_LOOP_4_1_mux1h_5_itm = MUX_v_40_12_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_1, attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_1,
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_1, attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_1,
      attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_1, attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_1,
      attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_1, attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_1,
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_1, attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_1,
      attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_1, {reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2});
  assign or_3156_nl = (fsm_output[6]) | (fsm_output[0]) | (~ (fsm_output[1]));
  assign or_3157_nl = (~ (fsm_output[6])) | (~ (fsm_output[0])) | (fsm_output[1]);
  assign mux_905_nl = MUX_s_1_2_2(or_3156_nl, or_3157_nl, fsm_output[7]);
  assign and_404_itm = (~(mux_905_nl | (fsm_output[8]))) & and_dcpl_364 & and_dcpl_194;
  assign rms_norm_16_variance_or_1_cse = and_dcpl_242 | (and_dcpl_239 & and_dcpl_182);
  assign nor_985_nl = ~((fsm_output[6]) | (fsm_output[3]) | (fsm_output[5]) | (fsm_output[0])
      | (fsm_output[1]) | (fsm_output[2]));
  assign and_1566_nl = (fsm_output[3]) & (fsm_output[5]) & (fsm_output[0]) & (fsm_output[1])
      & (~ (fsm_output[2]));
  assign nor_986_nl = ~((~ (fsm_output[3])) | (fsm_output[5]) | (fsm_output[0]) |
      (fsm_output[1]) | (~ (fsm_output[2])));
  assign mux_947_nl = MUX_s_1_2_2(and_1566_nl, nor_986_nl, fsm_output[6]);
  assign mux_948_nl = MUX_s_1_2_2(nor_985_nl, mux_947_nl, fsm_output[7]);
  assign GEMM_3D_FLOAT_LOOP_4_1_nand_itm = ~(mux_948_nl & and_dcpl_61);
  assign mux_941_nl = MUX_s_1_2_2(mux_tmp_916, or_1197_cse, fsm_output[4]);
  assign mux_939_nl = MUX_s_1_2_2(mux_tmp_936, or_1197_cse, fsm_output[4]);
  assign mux_940_nl = MUX_s_1_2_2(mux_939_nl, mux_tmp_937, or_1880_cse);
  assign mux_942_nl = MUX_s_1_2_2(mux_941_nl, mux_940_nl, fsm_output[0]);
  assign mux_938_nl = MUX_s_1_2_2(mux_tmp_937, mux_tmp_922, fsm_output[0]);
  assign mux_943_nl = MUX_s_1_2_2(mux_942_nl, mux_938_nl, fsm_output[1]);
  assign mux_933_nl = MUX_s_1_2_2(or_tmp_808, or_tmp_805, fsm_output[4]);
  assign mux_934_nl = MUX_s_1_2_2(mux_933_nl, mux_tmp_927, fsm_output[0]);
  assign mux_932_nl = MUX_s_1_2_2(or_tmp_805, or_tmp_812, fsm_output[4]);
  assign mux_935_nl = MUX_s_1_2_2(mux_934_nl, mux_932_nl, fsm_output[1]);
  assign mux_944_nl = MUX_s_1_2_2(mux_943_nl, mux_935_nl, fsm_output[5]);
  assign mux_928_nl = MUX_s_1_2_2(or_362_cse, or_361_cse, or_1879_cse);
  assign mux_929_nl = MUX_s_1_2_2(mux_928_nl, mux_tmp_927, fsm_output[0]);
  assign mux_930_nl = MUX_s_1_2_2(mux_tmp_915, mux_929_nl, fsm_output[1]);
  assign mux_931_nl = MUX_s_1_2_2(mux_tmp_908, mux_930_nl, fsm_output[5]);
  assign mux_945_nl = MUX_s_1_2_2(mux_944_nl, mux_931_nl, fsm_output[3]);
  assign mux_920_nl = MUX_s_1_2_2(mux_tmp_919, or_tmp_813, fsm_output[4]);
  assign mux_923_nl = MUX_s_1_2_2(mux_tmp_922, mux_920_nl, fsm_output[0]);
  assign mux_917_nl = MUX_s_1_2_2(mux_tmp_916, or_tmp_813, fsm_output[4]);
  assign mux_918_nl = MUX_s_1_2_2(mux_917_nl, mux_tmp_910, fsm_output[0]);
  assign mux_924_nl = MUX_s_1_2_2(mux_923_nl, mux_918_nl, fsm_output[1]);
  assign mux_925_nl = MUX_s_1_2_2(mux_924_nl, mux_tmp_915, fsm_output[5]);
  assign mux_912_nl = MUX_s_1_2_2(mux_tmp_908, mux_tmp_910, fsm_output[0]);
  assign mux_911_nl = MUX_s_1_2_2(mux_tmp_910, mux_tmp_908, fsm_output[0]);
  assign mux_913_nl = MUX_s_1_2_2(mux_912_nl, mux_911_nl, fsm_output[1]);
  assign mux_907_nl = MUX_s_1_2_2(mux_tmp_906, or_tmp_805, or_1867_cse);
  assign mux_914_nl = MUX_s_1_2_2(mux_913_nl, mux_907_nl, fsm_output[5]);
  assign mux_926_nl = MUX_s_1_2_2(mux_925_nl, mux_914_nl, fsm_output[3]);
  assign mux_946_nl = MUX_s_1_2_2(mux_945_nl, mux_926_nl, fsm_output[2]);
  assign GEMM_3D_FLOAT_LOOP_4_1_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & mux_946_nl;
  assign or_1907_cse = (fsm_output[2:1]!=2'b01);
  assign and_1572_cse = (fsm_output[2:0]==3'b111);
  assign or_1908_cse = (fsm_output[2:1]!=2'b00);
  assign and_1570_cse = (fsm_output[1]) & (fsm_output[2]) & (fsm_output[4]);
  assign nor_992_cse = ~((fsm_output[2]) | (fsm_output[4]));
  assign nand_240_cse = ~((fsm_output[1]) & (fsm_output[0]) & (fsm_output[2]) & (fsm_output[4]));
  assign mux_958_cse = MUX_s_1_2_2(or_tmp_48, or_133_cse, fsm_output[5]);
  assign or_1890_nl = (fsm_output[3]) | (fsm_output[5]) | (~ (fsm_output[0])) | (fsm_output[2])
      | (fsm_output[6]);
  assign or_3158_nl = (~ (fsm_output[2])) | (fsm_output[6]);
  assign nand_318_nl = ~((fsm_output[2]) & (fsm_output[6]));
  assign mux_950_nl = MUX_s_1_2_2(or_3158_nl, nand_318_nl, fsm_output[0]);
  assign or_1889_nl = (~ (fsm_output[3])) | (fsm_output[5]) | mux_950_nl;
  assign mux_951_nl = MUX_s_1_2_2(or_1890_nl, or_1889_nl, fsm_output[7]);
  assign nor_990_nl = ~((fsm_output[8]) | mux_951_nl);
  assign nor_988_nl = ~(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4 | (~ (fsm_output[0]))
      | (fsm_output[2]) | (fsm_output[6]));
  assign nor_989_nl = ~((fsm_output[0]) | (~ (fsm_output[2])) | (fsm_output[6]));
  assign mux_949_nl = MUX_s_1_2_2(nor_988_nl, nor_989_nl, fsm_output[5]);
  assign and_1568_nl = (~((~ (fsm_output[8])) | (fsm_output[7]) | (~ (fsm_output[3]))))
      & mux_949_nl;
  assign mux_952_nl = MUX_s_1_2_2(nor_990_nl, and_1568_nl, fsm_output[4]);
  assign and_416_itm = mux_952_nl & (fsm_output[1]);
  assign nand_47_nl = ~((fsm_output[5]) & nor_998_cse);
  assign mux_985_nl = MUX_s_1_2_2(nand_47_nl, or_tmp_798, fsm_output[3]);
  assign and_428_itm = (~ mux_985_nl) & and_dcpl_390;
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_cse = and_dcpl_382 | and_dcpl_386;
  assign or_3206_nl = (fsm_output[4:2]!=3'b110);
  assign or_3207_nl = (fsm_output[4:2]!=3'b001);
  assign mux_2236_nl = MUX_s_1_2_2(or_3206_nl, or_3207_nl, fsm_output[6]);
  assign nor_1314_cse = ~(mux_2236_nl | (fsm_output[8]));
  assign or_1923_nl = (fsm_output[3]) | (fsm_output[6]) | (fsm_output[8]);
  assign or_1922_nl = (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[8]));
  assign mux_978_nl = MUX_s_1_2_2(or_1923_nl, or_1922_nl, fsm_output[4]);
  assign or_1920_nl = (fsm_output[4]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[8]);
  assign mux_979_nl = MUX_s_1_2_2(mux_978_nl, or_1920_nl, fsm_output[2]);
  assign or_1919_nl = (~ (fsm_output[4])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (fsm_output[8]);
  assign or_1918_nl = (fsm_output[4]) | (~ (fsm_output[3])) | (~ (fsm_output[6]))
      | (fsm_output[8]);
  assign mux_977_nl = MUX_s_1_2_2(or_1919_nl, or_1918_nl, fsm_output[2]);
  assign mux_980_nl = MUX_s_1_2_2(mux_979_nl, mux_977_nl, fsm_output[7]);
  assign or_3159_nl = (fsm_output[1]) | mux_980_nl;
  assign or_1916_nl = (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[8]);
  assign nand_321_nl = ~(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4 & (fsm_output[3])
      & (~ (fsm_output[6])) & (fsm_output[8]));
  assign mux_976_nl = MUX_s_1_2_2(or_1916_nl, nand_321_nl, fsm_output[4]);
  assign or_3160_nl = (~ (fsm_output[1])) | (fsm_output[7]) | (fsm_output[2]) | mux_976_nl;
  assign mux_981_nl = MUX_s_1_2_2(or_3159_nl, or_3160_nl, fsm_output[0]);
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_5_itm = mux_981_nl | (fsm_output[5]);
  assign mux_969_nl = MUX_s_1_2_2(or_tmp_48, or_133_cse, and_1559_cse);
  assign mux_970_nl = MUX_s_1_2_2(mux_969_nl, mux_tmp_968, fsm_output[0]);
  assign nor_991_nl = ~(and_1570_cse | (fsm_output[8]));
  assign mux_971_nl = MUX_s_1_2_2(mux_970_nl, nor_991_nl, fsm_output[5]);
  assign mux_964_nl = MUX_s_1_2_2(and_dcpl_61, mux_528_cse, or_1908_cse);
  assign mux_963_nl = MUX_s_1_2_2(and_dcpl_61, mux_528_cse, or_1907_cse);
  assign mux_965_nl = MUX_s_1_2_2(mux_964_nl, mux_963_nl, fsm_output[0]);
  assign nand_319_nl = ~((~((fsm_output[1]) & (fsm_output[2]) & (fsm_output[4])))
      & (fsm_output[8]));
  assign mux_961_nl = MUX_s_1_2_2(mux_tmp_960, nand_319_nl, fsm_output[0]);
  assign mux_966_nl = MUX_s_1_2_2((~ mux_965_nl), mux_961_nl, fsm_output[5]);
  assign mux_972_nl = MUX_s_1_2_2(mux_971_nl, mux_966_nl, fsm_output[3]);
  assign or_1901_nl = nor_992_cse | (fsm_output[8]);
  assign or_1899_nl = and_1572_cse | (fsm_output[4]) | (fsm_output[8]);
  assign mux_957_nl = MUX_s_1_2_2(or_1901_nl, or_1899_nl, fsm_output[5]);
  assign mux_959_nl = MUX_s_1_2_2(mux_958_cse, mux_957_nl, fsm_output[3]);
  assign mux_973_nl = MUX_s_1_2_2(mux_972_nl, mux_959_nl, fsm_output[6]);
  assign or_1898_nl = (fsm_output[2]) | (fsm_output[4]) | (fsm_output[8]);
  assign mux_954_nl = MUX_s_1_2_2(or_1898_nl, or_tmp_833, or_1732_cse);
  assign mux_955_nl = MUX_s_1_2_2(or_tmp_757, mux_954_nl, fsm_output[5]);
  assign or_1895_nl = (fsm_output[5]) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_956_nl = MUX_s_1_2_2(mux_955_nl, or_1895_nl, fsm_output[3]);
  assign nand_46_nl = ~((fsm_output[6]) & (~ mux_956_nl));
  assign mux_974_nl = MUX_s_1_2_2(mux_973_nl, nand_46_nl, fsm_output[7]);
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & mux_974_nl;
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_7_cse = and_dcpl_328 & and_428_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_8_cse = and_dcpl_313 & and_428_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_9_cse = and_dcpl_587 & and_dcpl_190
      & and_428_itm;
  assign compute_sqrt_for_i_and_2_cse = (~ and_dcpl_557) & and_dcpl_414;
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c0 | and_dcpl_242 | LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c2
      | LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c3 | LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c5
      | and_dcpl_410 | LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c7 | and_dcpl_414);
  assign compute_sqrt_for_i_and_cse = and_dcpl_201 & and_1474_cse & and_dcpl_199
      & LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c7;
  assign nor_1311_nl = ~((fsm_output[1:0]!=2'b00) | or_dcpl_1050);
  assign mux_2227_nl = MUX_s_1_2_2(nor_1311_nl, mux_tmp_1451, fsm_output[5]);
  assign mux_2228_nl = MUX_s_1_2_2(mux_2227_nl, and_tmp_42, fsm_output[3]);
  assign mux_2229_nl = MUX_s_1_2_2(mux_2228_nl, (~ or_tmp_755), fsm_output[6]);
  assign compute_sqrt_for_i_and_4_cse = mux_2229_nl & and_dcpl_295 & LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c7;
  assign compute_sqrt_for_i_and_5_cse = (and_dcpl_328 | and_dcpl_635) & LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c7;
  assign and_1773_cse = (fsm_output[3:2]==2'b11);
  assign or_1983_cse = (fsm_output[7:6]!=2'b01);
  assign or_1985_cse = (fsm_output[7:5]!=3'b011);
  assign or_1984_cse = (fsm_output[7:6]!=2'b00);
  assign nor_1026_cse = ~((fsm_output[0]) | (fsm_output[5]));
  assign for_for_and_13_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 &
      (and_dcpl_415 | for_for_strm_in_tmp_sva_31_2_mx0c1);
  assign and_474_rgt = and_dcpl_342 & and_dcpl_336 & and_dcpl_433;
  assign and_476_rgt = or_dcpl_1071 & and_dcpl_185 & and_dcpl_422;
  assign and_480_rgt = and_dcpl_350 & and_dcpl_190;
  assign for_for_and_14_rgt = (~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd | reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1))
      & and_dcpl_442;
  assign for_for_and_15_rgt = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd)
      & and_dcpl_442;
  assign for_for_and_16_rgt = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1)
      & and_dcpl_442;
  assign for_for_and_17_rgt = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      & and_dcpl_442;
  assign and_485_rgt = and_dcpl_241 & (fsm_output[5]) & SOFTMAX_LOOP_3_acc_3_itm_40_1
      & (fsm_output[3]) & and_dcpl_45;
  assign and_486_rgt = and_dcpl_376 & and_dcpl_221;
  assign for_for_or_1_rgt = and_dcpl_448 | (and_dcpl_449 & and_dcpl_200 & and_dcpl_261);
  assign nand_328_nl = ~((fsm_output[2]) & (fsm_output[5]) & (fsm_output[3]) & (fsm_output[7]));
  assign or_2016_nl = (fsm_output[5]) | (fsm_output[3]) | (fsm_output[7]);
  assign or_2015_nl = SOFTMAX_LOOP_3_acc_3_itm_40_1 | not_tmp_549;
  assign mux_1068_nl = MUX_s_1_2_2(or_2016_nl, or_2015_nl, fsm_output[0]);
  assign or_2014_nl = (fsm_output[0]) | not_tmp_549;
  assign mux_1069_nl = MUX_s_1_2_2(mux_1068_nl, or_2014_nl, fsm_output[2]);
  assign mux_1070_nl = MUX_s_1_2_2(nand_328_nl, mux_1069_nl, fsm_output[1]);
  assign or_2013_nl = (~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 | reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1))
      | (~ (fsm_output[0])) | (fsm_output[5]) | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1066_nl = MUX_s_1_2_2(or_2013_nl, or_tmp_938, fsm_output[2]);
  assign or_2007_nl = (fsm_output[3]) | (~ (fsm_output[7]));
  assign or_2006_nl = (fsm_output[3]) | (fsm_output[7]);
  assign mux_1064_nl = MUX_s_1_2_2(or_2007_nl, or_2006_nl, fsm_output[5]);
  assign or_2008_nl = (fsm_output[0]) | mux_1064_nl;
  assign mux_1065_nl = MUX_s_1_2_2(or_tmp_938, or_2008_nl, fsm_output[2]);
  assign mux_1067_nl = MUX_s_1_2_2(mux_1066_nl, mux_1065_nl, fsm_output[1]);
  assign mux_1071_nl = MUX_s_1_2_2(mux_1070_nl, mux_1067_nl, fsm_output[4]);
  assign nand_329_nl = ~((fsm_output[4]) & (~ (fsm_output[1])) & (fsm_output[2])
      & (fsm_output[0]) & (fsm_output[5]) & (~ (fsm_output[3])) & (fsm_output[7]));
  assign mux_1072_nl = MUX_s_1_2_2(mux_1071_nl, nand_329_nl, fsm_output[6]);
  assign QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (mux_1072_nl | (fsm_output[8]));
  assign and_37_cse = (RMS_NORM_LOOP_2_2_i_4_0_sva_1[4]) & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  assign GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_8_seb = ~(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva_mx0w3
      & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  assign mux_1114_nl = MUX_s_1_2_2((~ nor_tmp_289), mux_tmp_1113, fsm_output[0]);
  assign mux_1115_nl = MUX_s_1_2_2(mux_1114_nl, or_tmp_992, fsm_output[6]);
  assign mux_1116_nl = MUX_s_1_2_2(or_tmp_993, mux_1115_nl, fsm_output[7]);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_and_37_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~ or_dcpl_1068) | apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c0
      | apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c1 | and_dcpl_477 | and_dcpl_220
      | and_dcpl_222 | and_dcpl_187) & (~((~ mux_1116_nl) & and_dcpl_478));
  assign or_2081_nl = (fsm_output[1]) | or_dcpl_1050;
  assign or_2080_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (~ (fsm_output[4]));
  assign mux_1117_nl = MUX_s_1_2_2(or_2081_nl, or_2080_nl, fsm_output[0]);
  assign mux_1118_nl = MUX_s_1_2_2(mux_1117_nl, or_tmp_992, fsm_output[6]);
  assign mux_1119_nl = MUX_s_1_2_2(or_tmp_993, mux_1118_nl, fsm_output[7]);
  assign attention_2_1_16_16_4_4_attn_output_and_25_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~((~ mux_1119_nl) & and_dcpl_478));
  assign or_3212_tmp = (and_dcpl_1233 & GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva_mx0w0)
      | mux_tmp_1163;
  assign or_3213_tmp = (and_dcpl_1233 & GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva_mx0w0)
      | mux_tmp_1163;
  assign or_3214_tmp = (and_dcpl_1233 & GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva_mx0w0)
      | attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c10;
  assign nor_366_cse = ~((fsm_output[1:0]!=2'b10));
  assign or_3167_cse = (fsm_output[2:1]!=2'b10);
  assign or_2154_cse = (~ (fsm_output[5])) | (fsm_output[7]);
  assign nor_1044_cse = ~((~ (fsm_output[3])) | (~ (fsm_output[1])) | (~ (fsm_output[2]))
      | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1045_cse = ~((~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[1])
      | (~ (fsm_output[2])) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1208_nl = MUX_s_1_2_2(and_dcpl_449, and_dcpl_263, fsm_output[1]);
  assign mux_1209_nl = MUX_s_1_2_2(and_dcpl_341, mux_1208_nl, fsm_output[3]);
  assign mux_1210_nl = MUX_s_1_2_2(mux_1209_nl, nor_1044_cse, fsm_output[6]);
  assign mux_1211_nl = MUX_s_1_2_2(mux_1210_nl, nor_1045_cse, fsm_output[7]);
  assign and_581_ssc = mux_1211_nl & and_dcpl_338;
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_nand_seb = ~(and_dcpl_381 & nor_777_cse
      & and_dcpl_198);
  assign nor_1046_nl = ~((fsm_output[6]) | (fsm_output[0]) | (fsm_output[1]) | (~
      (fsm_output[2])));
  assign and_1597_nl = (fsm_output[6]) & (fsm_output[0]) & (fsm_output[1]) & (~ (fsm_output[2]));
  assign mux_1212_nl = MUX_s_1_2_2(nor_1046_nl, and_1597_nl, fsm_output[7]);
  assign and_585_seb = mux_1212_nl & and_dcpl_201 & and_dcpl_189;
  assign mux_1231_nl = MUX_s_1_2_2(mux_tmp_1229, mux_tmp_1219, fsm_output[1]);
  assign mux_1230_nl = MUX_s_1_2_2(mux_tmp_1229, mux_tmp_1219, fsm_output[2]);
  assign mux_1232_nl = MUX_s_1_2_2(mux_1231_nl, mux_1230_nl, fsm_output[0]);
  assign mux_1233_nl = MUX_s_1_2_2(mux_1232_nl, or_1795_cse, fsm_output[6]);
  assign mux_1226_nl = MUX_s_1_2_2(mux_tmp_1218, or_tmp_1051, fsm_output[2]);
  assign mux_1225_nl = MUX_s_1_2_2(mux_tmp_1218, or_2154_cse, fsm_output[2]);
  assign mux_1227_nl = MUX_s_1_2_2(mux_1226_nl, mux_1225_nl, or_1732_cse);
  assign or_2152_nl = (~((fsm_output[2]) | (~ (fsm_output[7])))) | (fsm_output[8]);
  assign or_2151_nl = (~((fsm_output[2]) | (~ (fsm_output[5])) | (~ (fsm_output[7]))))
      | (fsm_output[8]);
  assign mux_1223_nl = MUX_s_1_2_2(or_2152_nl, or_2151_nl, fsm_output[1]);
  assign or_2150_nl = (or_3167_cse & (fsm_output[5]) & (fsm_output[7])) | (fsm_output[8]);
  assign mux_1224_nl = MUX_s_1_2_2(mux_1223_nl, or_2150_nl, fsm_output[0]);
  assign mux_1228_nl = MUX_s_1_2_2(mux_1227_nl, mux_1224_nl, fsm_output[6]);
  assign mux_1234_nl = MUX_s_1_2_2(mux_1233_nl, mux_1228_nl, fsm_output[4]);
  assign mux_1220_nl = MUX_s_1_2_2(mux_tmp_1219, mux_tmp_1218, and_1559_cse);
  assign or_2145_nl = (~ (fsm_output[2])) | (fsm_output[5]);
  assign mux_1216_nl = MUX_s_1_2_2(or_361_cse, or_362_cse, or_2145_nl);
  assign mux_1217_nl = MUX_s_1_2_2(or_1795_cse, mux_1216_nl, nor_366_cse);
  assign mux_1221_nl = MUX_s_1_2_2(mux_1220_nl, mux_1217_nl, fsm_output[6]);
  assign or_2142_nl = (fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[8]));
  assign mux_1213_nl = MUX_s_1_2_2(or_tmp_1051, or_2142_nl, fsm_output[1]);
  assign or_2140_nl = and_1559_cse | (~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[8]));
  assign mux_1214_nl = MUX_s_1_2_2(mux_1213_nl, or_2140_nl, fsm_output[0]);
  assign or_2138_nl = ((fsm_output[5]) & (fsm_output[7])) | (fsm_output[8]);
  assign mux_1215_nl = MUX_s_1_2_2(mux_1214_nl, or_2138_nl, fsm_output[6]);
  assign mux_1222_nl = MUX_s_1_2_2(mux_1221_nl, mux_1215_nl, fsm_output[4]);
  assign mux_1235_nl = MUX_s_1_2_2(mux_1234_nl, mux_1222_nl, fsm_output[3]);
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_1_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & mux_1235_nl;
  assign attention_abs_qelse_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~(((and_1637_cse | (fsm_output[3])) ^ (fsm_output[4])) & and_dcpl_270));
  assign compute_sqrt_guess_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((and_dcpl_192 & and_dcpl_209) | and_dcpl_290);
  assign nor_1229_cse = ~(reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign and_1191_rgt = and_dcpl_1061 & and_dcpl_45 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      & nor_1229_cse & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd;
  assign mux_1310_nl = MUX_s_1_2_2(or_tmp_611, or_tmp_1128, fsm_output[3]);
  assign and_622_rgt = (~ mux_1310_nl) & and_dcpl_581;
  assign operator_40_24_true_AC_TRN_AC_WRAP_1_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~(or_dcpl_1040 & and_dcpl_191 & and_dcpl_321 & and_dcpl_1141));
  assign operator_40_24_true_AC_TRN_AC_WRAP_1_conc_1_itm_11_0 = MUX_v_12_16_2(12'b011110001010,
      12'b011101010010, 12'b100000010100, 12'b011100010010, 12'b011100110010, 12'b100000011110,
      12'b011101100011, 12'b100000101100, 12'b011111110100, 12'b011100010000, 12'b011110000101,
      12'b100001110110, 12'b011101111110, 12'b011110001010, 12'b100000111010, 12'b100001001110,
      {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
  assign operator_40_24_true_AC_TRN_AC_WRAP_1_conc_3_itm_8_0 = MUX_v_9_16_2(9'b011001100,
      9'b001101100, 9'b101011100, 9'b100110000, 9'b010100011, 9'b101100000, 9'b011001100,
      9'b101000111, 9'b110000011, 9'b010111100, 9'b010001100, 9'b100000000, 9'b011000000,
      9'b000100111, 9'b110111000, 9'b101110011, {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
      , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
  assign or_3174_nl = (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign nand_344_nl = ~((fsm_output[6]) & (fsm_output[3]) & (fsm_output[2]));
  assign mux_1308_nl = MUX_s_1_2_2(or_3174_nl, nand_344_nl, fsm_output[7]);
  assign and_615_itm = (~(mux_1308_nl | (fsm_output[8]))) & and_1651_cse & nor_1026_cse;
  assign operator_40_24_true_AC_TRN_AC_WRAP_1_and_4_cse = (~ and_1191_rgt) & and_622_rgt;
  assign attention_2_1_16_16_4_4_quantized_hidden_states_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1087 | and_dcpl_618)) | or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_cse = QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1
      & and_dcpl_619;
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_cse = (~
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1) & and_dcpl_619;
  assign attention_2_1_16_16_4_4_quantized_hidden_states_and_1_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1086 | and_dcpl_618)) | or_dcpl_1104);
  assign attention_2_1_16_16_4_4_quantized_hidden_states_and_2_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1067 | and_dcpl_618)) | or_dcpl_1104);
  assign attention_2_1_16_16_4_4_quantized_hidden_states_and_3_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1079 | and_dcpl_618)) | or_dcpl_1104);
  assign or_3185_cse = (fsm_output[2:0]!=3'b000);
  assign and_1637_cse = or_1732_cse & (fsm_output[2]);
  assign RMS_NORM_LOOP_2_2_i_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (and_dcpl_477 | RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c1 | and_dcpl_410 | and_dcpl_620
      | RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c4 | and_dcpl_255);
  assign RMS_NORM_LOOP_2_2_i_and_9_cse = and_dcpl_564 & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1)
      & and_dcpl_620;
  assign or_2249_cse = (fsm_output[7:6]!=2'b10);
  assign and_633_itm = and_dcpl_588 & and_dcpl_592;
  assign and_654_itm = and_dcpl_588 & and_dcpl_613;
  assign and_648_itm = and_dcpl_588 & and_dcpl_607;
  assign and_642_itm = and_dcpl_588 & and_dcpl_601;
  assign and_636_itm = and_dcpl_588 & and_dcpl_595;
  assign and_629_itm = and_dcpl_588 & and_dcpl_586;
  assign and_639_itm = and_dcpl_588 & and_dcpl_598;
  assign and_645_itm = and_dcpl_588 & and_dcpl_604;
  assign and_651_itm = and_dcpl_588 & and_dcpl_610;
  assign and_657_itm = and_dcpl_588 & and_dcpl_616;
  assign and_1638_cse = (fsm_output[3:1]==3'b111);
  assign nor_1106_cse = ~((fsm_output[2:0]!=3'b000));
  assign and_937_ssc = (~(mux_tmp_1426 | (fsm_output[8]))) & and_dcpl_338 & and_dcpl_45;
  assign nand_71_nl = ~((fsm_output[6]) & (fsm_output[3]) & (~(and_1474_cse | (~
      (fsm_output[2])) | (fsm_output[4]))));
  assign mux_1636_nl = MUX_s_1_2_2(or_tmp_1221, or_tmp_1128, fsm_output[0]);
  assign mux_1637_nl = MUX_s_1_2_2(or_tmp_1203, mux_1636_nl, fsm_output[3]);
  assign or_2563_nl = (fsm_output[6]) | mux_1637_nl;
  assign mux_1638_nl = MUX_s_1_2_2(nand_71_nl, or_2563_nl, fsm_output[7]);
  assign nor_1324_seb = ~(mux_1638_nl | or_1851_cse);
  assign and_679_nl = (fsm_output[5]) & mux_tmp_1451;
  assign mux_1452_nl = MUX_s_1_2_2(and_679_nl, and_tmp_42, fsm_output[3]);
  assign mux_1453_nl = MUX_s_1_2_2(mux_1452_nl, (~ or_tmp_755), fsm_output[6]);
  assign CACHE_UPDATE_LOOP_3_k_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~(mux_1453_nl & and_dcpl_295));
  assign QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_or_cse = and_dcpl_888
      | (and_dcpl_362 & and_dcpl_237);
  assign nand_197_cse = ~((fsm_output[1:0]==2'b11));
  assign nor_777_cse = ~((fsm_output[1:0]!=2'b00));
  assign nand_350_nl = ~(or_2500_cse & (fsm_output[7]));
  assign or_2355_nl = (fsm_output[1]) | (~ (fsm_output[7]));
  assign mux_1456_nl = MUX_s_1_2_2(nand_350_nl, or_2355_nl, fsm_output[0]);
  assign nor_1115_nl = ~((fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | mux_1456_nl);
  assign nor_1116_nl = ~((~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[0])
      | (fsm_output[1]) | (fsm_output[7]));
  assign nor_1114_nl = ~(nor_777_cse | (fsm_output[7]));
  assign mux_1454_nl = MUX_s_1_2_2(nor_1114_nl, (fsm_output[7]), fsm_output[6]);
  assign nor_1117_nl = ~((fsm_output[3]) | (~ mux_1454_nl));
  assign mux_1455_nl = MUX_s_1_2_2(nor_1116_nl, nor_1117_nl, fsm_output[2]);
  assign mux_1457_nl = MUX_s_1_2_2(nor_1115_nl, mux_1455_nl, fsm_output[5]);
  assign GEMM_3D_FLOAT_LOOP_1_i_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((mux_1457_nl & and_dcpl_201) | GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c1
      | GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c2);
  assign nand_126_nl = ~((fsm_output[5:3]==3'b111));
  assign mux_1490_nl = MUX_s_1_2_2(nand_126_nl, mux_tmp_1489, fsm_output[6]);
  assign input_and_28_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~((~
      mux_1490_nl) & and_dcpl_26));
  assign and_699_ssc = or_dcpl_1116 & and_dcpl_202 & and_dcpl_642;
  assign and_745_ssc = or_dcpl_1131 & and_dcpl_202 & and_dcpl_642;
  assign or_2456_cse = (fsm_output[6]) | (~ (fsm_output[8]));
  assign or_2457_cse = (fsm_output[8:6]!=3'b001);
  assign or_2455_cse = (fsm_output[6]) | (fsm_output[8]);
  assign or_2460_cse = (fsm_output[4]) | (~ (fsm_output[7])) | (~ (fsm_output[6]))
      | (fsm_output[8]);
  assign or_2451_cse = (fsm_output[4]) | (~ (fsm_output[7])) | (fsm_output[6]) |
      (fsm_output[8]);
  assign mux_1522_cse = MUX_s_1_2_2(or_2456_cse, or_2455_cse, fsm_output[7]);
  assign or_2443_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[4]);
  assign mux_1513_cse = MUX_s_1_2_2(or_2443_nl, or_tmp_1128, fsm_output[0]);
  assign mux_1496_nl = MUX_s_1_2_2(or_tmp_931, or_2154_cse, fsm_output[4]);
  assign or_2429_nl = (fsm_output[6]) | mux_1496_nl;
  assign or_2426_nl = (fsm_output[2]) | (~ (fsm_output[3])) | (fsm_output[0]);
  assign mux_1497_nl = MUX_s_1_2_2(or_2429_nl, or_tmp_1291, or_2426_nl);
  assign nand_354_nl = ~((fsm_output[4]) & (fsm_output[5]) & (fsm_output[7]));
  assign mux_1492_nl = MUX_s_1_2_2(or_tmp_930, nand_354_nl, fsm_output[6]);
  assign mux_1493_nl = MUX_s_1_2_2(or_tmp_1291, mux_1492_nl, fsm_output[0]);
  assign nand_355_nl = ~((fsm_output[7:4]==4'b0111));
  assign mux_1494_nl = MUX_s_1_2_2(mux_1493_nl, nand_355_nl, fsm_output[3]);
  assign mux_1495_nl = MUX_s_1_2_2(or_tmp_1291, mux_1494_nl, fsm_output[2]);
  assign mux_1498_nl = MUX_s_1_2_2(mux_1497_nl, mux_1495_nl, fsm_output[1]);
  assign nor_1138_m1c = ~(mux_1498_nl | (fsm_output[8]));
  assign or_2442_nl = (fsm_output[3:2]!=2'b00) | (~ RESHAPE_2D_TO_3D_LOOP_2_2_and_cse)
      | (~ (fsm_output[4])) | (~ (fsm_output[7])) | (fsm_output[6]) | (fsm_output[8]);
  assign mux_1510_nl = MUX_s_1_2_2(or_2442_nl, or_tmp_1296, fsm_output[5]);
  assign or_2441_nl = (~ RESHAPE_2D_TO_3D_LOOP_2_2_and_cse) | (~ (fsm_output[4]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (fsm_output[8]);
  assign mux_1507_nl = MUX_s_1_2_2(or_2441_nl, mux_tmp_1519, fsm_output[3]);
  assign or_2438_nl = (~ (z_out_4[2])) | (~ (fsm_output[4])) | (~ (fsm_output[7]))
      | (fsm_output[6]) | (fsm_output[8]);
  assign mux_1505_nl = MUX_s_1_2_2(or_2438_nl, or_2451_cse, fsm_output[3]);
  assign mux_1508_nl = MUX_s_1_2_2(mux_1507_nl, mux_1505_nl, fsm_output[2]);
  assign or_2436_nl = reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 | (fsm_output[8:6]!=3'b010);
  assign mux_1503_nl = MUX_s_1_2_2(or_2436_nl, or_1197_cse, fsm_output[4]);
  assign mux_1504_nl = MUX_s_1_2_2(or_2451_cse, mux_1503_nl, fsm_output[3]);
  assign nand_64_nl = ~((fsm_output[2]) & (~ mux_1504_nl));
  assign mux_1509_nl = MUX_s_1_2_2(mux_1508_nl, nand_64_nl, fsm_output[5]);
  assign mux_1511_nl = MUX_s_1_2_2(mux_1510_nl, mux_1509_nl, fsm_output[1]);
  assign mux_1500_nl = MUX_s_1_2_2(or_2460_cse, mux_2092_cse, fsm_output[3]);
  assign or_2431_nl = (~ (fsm_output[3])) | (~ (fsm_output[4])) | (~ (fsm_output[7]))
      | (fsm_output[6]) | (fsm_output[8]);
  assign mux_1501_nl = MUX_s_1_2_2(mux_1500_nl, or_2431_nl, fsm_output[2]);
  assign mux_1502_nl = MUX_s_1_2_2(mux_1501_nl, or_tmp_1296, fsm_output[5]);
  assign nand_63_nl = ~((fsm_output[1]) & (~ mux_1502_nl));
  assign mux_1512_itm = MUX_s_1_2_2(mux_1511_nl, nand_63_nl, fsm_output[0]);
  assign mux_1529_nl = MUX_s_1_2_2(or_2460_cse, mux_tmp_1519, fsm_output[3]);
  assign or_2459_nl = (fsm_output[3]) | mux_tmp_1519;
  assign mux_1530_nl = MUX_s_1_2_2(mux_1529_nl, or_2459_nl, fsm_output[0]);
  assign or_2458_nl = (~ (fsm_output[4])) | (~ (fsm_output[7])) | (fsm_output[6])
      | (fsm_output[8]);
  assign mux_1527_nl = MUX_s_1_2_2(or_2458_nl, mux_tmp_1519, fsm_output[3]);
  assign mux_1528_nl = MUX_s_1_2_2(or_tmp_1320, mux_1527_nl, fsm_output[0]);
  assign mux_1531_nl = MUX_s_1_2_2(mux_1530_nl, mux_1528_nl, fsm_output[1]);
  assign mux_1532_nl = MUX_s_1_2_2(mux_1531_nl, or_tmp_1316, fsm_output[5]);
  assign mux_1523_nl = MUX_s_1_2_2(or_2457_cse, mux_1522_cse, fsm_output[4]);
  assign mux_1524_nl = MUX_s_1_2_2(mux_tmp_1519, mux_1523_nl, fsm_output[3]);
  assign mux_1520_nl = MUX_s_1_2_2(mux_tmp_1519, or_2451_cse, fsm_output[3]);
  assign mux_1521_nl = MUX_s_1_2_2(or_tmp_1320, mux_1520_nl, fsm_output[0]);
  assign mux_1525_nl = MUX_s_1_2_2(mux_1524_nl, mux_1521_nl, fsm_output[1]);
  assign or_2448_nl = (~((fsm_output[4:3]!=2'b00))) | (fsm_output[8:6]!=3'b010);
  assign mux_1517_nl = MUX_s_1_2_2(or_tmp_1316, or_2448_nl, fsm_output[0]);
  assign or_2446_nl = (~((~((fsm_output[0]) | (~ reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1)
      | (~ (fsm_output[3])))) | (fsm_output[4]))) | (fsm_output[8:6]!=3'b010);
  assign mux_1518_nl = MUX_s_1_2_2(mux_1517_nl, or_2446_nl, fsm_output[1]);
  assign mux_1526_nl = MUX_s_1_2_2(mux_1525_nl, mux_1518_nl, fsm_output[5]);
  assign mux_1533_nl = MUX_s_1_2_2(mux_1532_nl, mux_1526_nl, fsm_output[2]);
  assign APPLY_ROTARY_POS_EMB_LOOP_1_i_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & mux_1533_nl;
  assign mux_1540_nl = MUX_s_1_2_2(not_tmp_699, or_tmp_1132, fsm_output[7]);
  assign mux_1539_nl = MUX_s_1_2_2(not_tmp_699, or_tmp_1218, fsm_output[7]);
  assign mux_1541_nl = MUX_s_1_2_2(mux_1540_nl, mux_1539_nl, reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign nor_1144_itm = ~(mux_1541_nl | (fsm_output[8]));
  assign attention_2_1_16_16_4_4_q_proj_and_4_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((and_dcpl_588 & and_dcpl_721) | and_dcpl_240 | and_dcpl_626);
  assign attention_2_1_16_16_4_4_v_proj_re_and_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (and_dcpl_619 | and_dcpl_725 | and_dcpl_726 | and_dcpl_410);
  assign and_1651_cse = (fsm_output[4]) & (fsm_output[1]);
  assign or_2480_cse = (fsm_output[4]) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[8]);
  assign mux_1551_cse = MUX_s_1_2_2(or_tmp_464, or_2456_cse, fsm_output[5]);
  assign or_2481_cse = and_1651_cse | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[8]);
  assign mux_1559_cse = MUX_s_1_2_2(nand_tmp_66, mux_tmp_1549, fsm_output[4]);
  assign mux_1557_cse = MUX_s_1_2_2(mux_tmp_1549, mux_tmp_1548, and_1651_cse);
  assign and_1652_nl = (fsm_output[1]) & (fsm_output[5]);
  assign mux_1554_nl = MUX_s_1_2_2(mux_tmp_121, or_tmp_464, and_1652_nl);
  assign mux_1555_cse = MUX_s_1_2_2(mux_tmp_1549, mux_1554_nl, fsm_output[4]);
  assign mux_1552_nl = MUX_s_1_2_2(nand_tmp_66, mux_1551_cse, fsm_output[1]);
  assign mux_1550_nl = MUX_s_1_2_2(mux_tmp_1549, mux_tmp_1548, fsm_output[1]);
  assign mux_1553_cse = MUX_s_1_2_2(mux_1552_nl, mux_1550_nl, fsm_output[4]);
  assign or_2479_nl = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[0]);
  assign mux_1546_cse = MUX_s_1_2_2(or_2481_cse, or_2480_cse, or_2479_nl);
  assign mux_1564_nl = MUX_s_1_2_2(or_tmp_611, or_tmp_330, fsm_output[3]);
  assign attention_2_1_16_16_4_4_q_proj_re_and_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~((~ mux_1564_nl) & and_dcpl_581));
  assign or_2486_cse = reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd!=3'b100);
  assign or_2493_nl = (fsm_output[5]) | nor_tmp_285;
  assign mux_1580_nl = MUX_s_1_2_2(or_2493_nl, or_2699_cse, fsm_output[3]);
  assign or_2494_nl = (fsm_output[6]) | mux_1580_nl;
  assign mux_1581_nl = MUX_s_1_2_2(not_tmp_253, or_2494_nl, fsm_output[7]);
  assign attention_2_1_16_16_4_4_k_proj_re_and_1_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (mux_1581_nl | (fsm_output[8]));
  assign nand_381_cse = ~((fsm_output[4:3]==2'b11));
  assign or_3039_cse = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b00)
      | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  assign APPLY_ROTARY_POS_EMB_LOOP_6_k_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c0 | and_dcpl_726 | APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c2
      | APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c3 | APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c4);
  assign nand_365_cse = ~((fsm_output[7]) & (~(((RESHAPE_2D_TO_3D_LOOP_2_2_and_cse
      | (fsm_output[3:0]!=4'b0000)) & (fsm_output[4])) | (fsm_output[5]))));
  assign or_2566_nl = (fsm_output[5:4]!=2'b10);
  assign mux_1639_cse = MUX_s_1_2_2(or_2699_cse, or_2566_nl, fsm_output[1]);
  assign or_2576_nl = RESHAPE_2D_TO_3D_LOOP_2_2_and_cse | (fsm_output[2]) | (fsm_output[3])
      | (fsm_output[0]);
  assign mux_1645_cse = MUX_s_1_2_2(or_2481_cse, or_2480_cse, or_2576_nl);
  assign mux_1811_nl = MUX_s_1_2_2(mux_806_cse, or_1983_cse, fsm_output[1]);
  assign mux_1810_nl = MUX_s_1_2_2(or_2249_cse, mux_806_cse, fsm_output[1]);
  assign mux_1812_cse = MUX_s_1_2_2(mux_1811_nl, mux_1810_nl, fsm_output[0]);
  assign or_2638_nl = (fsm_output[3:0]!=4'b0000);
  assign mux_1809_cse = MUX_s_1_2_2(mux_806_cse, or_1983_cse, or_2638_nl);
  assign or_2671_cse = (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b01) | reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1
      | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]);
  assign or_2699_cse = (fsm_output[5:4]!=2'b00);
  assign and_1034_itm = and_dcpl_732 & and_dcpl_987;
  assign mux_1964_nl = MUX_s_1_2_2(mux_1559_cse, mux_1557_cse, and_1773_cse);
  assign mux_1959_nl = MUX_s_1_2_2(or_tmp_464, mux_tmp_121, or_2699_cse);
  assign mux_1958_nl = MUX_s_1_2_2(mux_tmp_1549, mux_tmp_1548, fsm_output[4]);
  assign mux_1960_nl = MUX_s_1_2_2(mux_1959_nl, mux_1958_nl, fsm_output[1]);
  assign mux_1954_nl = MUX_s_1_2_2(mux_1551_cse, mux_tmp_1548, fsm_output[4]);
  assign mux_1957_nl = MUX_s_1_2_2(mux_1559_cse, mux_1954_nl, fsm_output[1]);
  assign nor_540_nl = ~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b10));
  assign mux_1961_nl = MUX_s_1_2_2(mux_1960_nl, mux_1957_nl, nor_540_nl);
  assign mux_1962_nl = MUX_s_1_2_2(mux_1559_cse, mux_1961_nl, and_1773_cse);
  assign mux_1965_nl = MUX_s_1_2_2(mux_1964_nl, mux_1962_nl, fsm_output[0]);
  assign or_2696_nl = ((fsm_output[4:3]==2'b11)) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[8]);
  assign or_2695_nl = (~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 | reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      | (fsm_output[1]) | (~ (fsm_output[4])))) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[8]);
  assign mux_1948_nl = MUX_s_1_2_2(or_2695_nl, or_2481_cse, fsm_output[2]);
  assign mux_1949_nl = MUX_s_1_2_2(mux_1948_nl, or_2480_cse, fsm_output[3]);
  assign mux_1950_nl = MUX_s_1_2_2(or_2696_nl, mux_1949_nl, fsm_output[0]);
  assign mux_1966_itm = MUX_s_1_2_2(mux_1965_nl, mux_1950_nl, fsm_output[7]);
  assign and_1037_itm = and_dcpl_743 & and_dcpl_551 & and_dcpl_825;
  assign and_1042_ssc = and_dcpl_732 & and_dcpl_57 & (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[1]))
      & and_dcpl_651;
  assign nor_551_nl = ~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b00) | reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1
      | (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0])));
  assign mux_1982_nl = MUX_s_1_2_2(mux_806_cse, mux_1812_cse, nor_551_nl);
  assign mux_1983_nl = MUX_s_1_2_2(or_2249_cse, mux_1982_nl, and_1773_cse);
  assign or_2712_nl = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 | reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      | (fsm_output[1:0]!=2'b01);
  assign mux_1976_nl = MUX_s_1_2_2(or_1983_cse, mux_806_cse, or_2712_nl);
  assign mux_1975_nl = MUX_s_1_2_2(mux_806_cse, or_1983_cse, and_1474_cse);
  assign mux_1977_nl = MUX_s_1_2_2(mux_1976_nl, mux_1975_nl, fsm_output[2]);
  assign mux_1978_nl = MUX_s_1_2_2(mux_1977_nl, or_1983_cse, fsm_output[3]);
  assign mux_1984_nl = MUX_s_1_2_2(mux_1983_nl, mux_1978_nl, fsm_output[4]);
  assign mux_1985_nl = MUX_s_1_2_2(mux_1984_nl, or_1983_cse, fsm_output[5]);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_and_16_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (mux_1985_nl | (fsm_output[8]));
  assign or_2717_cse = (fsm_output[5]) | mux_806_cse;
  assign mux_1995_nl = MUX_s_1_2_2(mux_tmp_1993, mux_tmp_1990, fsm_output[2]);
  assign mux_1994_nl = MUX_s_1_2_2(mux_tmp_1993, or_2717_cse, and_1559_cse);
  assign nor_552_nl = ~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b11) | (~ (fsm_output[0])));
  assign mux_1996_nl = MUX_s_1_2_2(mux_1995_nl, mux_1994_nl, nor_552_nl);
  assign mux_1997_nl = MUX_s_1_2_2(mux_tmp_1993, mux_1996_nl, fsm_output[3]);
  assign or_2716_nl = (~ (fsm_output[1])) | (fsm_output[5]);
  assign mux_1988_nl = MUX_s_1_2_2(mux_806_cse, or_1983_cse, or_2716_nl);
  assign or_2715_nl = (fsm_output[1]) | (fsm_output[5]);
  assign mux_1987_nl = MUX_s_1_2_2(mux_806_cse, or_1983_cse, or_2715_nl);
  assign mux_1989_nl = MUX_s_1_2_2(mux_1988_nl, mux_1987_nl, fsm_output[2]);
  assign mux_1991_nl = MUX_s_1_2_2(mux_tmp_1990, mux_1989_nl, fsm_output[0]);
  assign mux_1992_nl = MUX_s_1_2_2(mux_1991_nl, or_1983_cse, fsm_output[3]);
  assign mux_1998_nl = MUX_s_1_2_2(mux_1997_nl, mux_1992_nl, fsm_output[4]);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_and_17_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1068 | (~(mux_1998_nl | (fsm_output[8]))))) | and_dcpl_619 |
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1 | and_dcpl_1003);
  assign and_1762_cse = (fsm_output[5:4]==2'b11);
  assign or_2742_cse = (~ (fsm_output[4])) | (~ (fsm_output[6])) | (fsm_output[8]);
  assign or_2736_cse = (fsm_output[4]) | (fsm_output[6]) | (~ (fsm_output[8]));
  assign or_2739_cse = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b01);
  assign mux_2024_cse = MUX_s_1_2_2(or_tmp_464, mux_tmp_121, fsm_output[4]);
  assign mux_2025_cse = MUX_s_1_2_2(mux_2024_cse, or_2736_cse, fsm_output[5]);
  assign mux_2032_cse = MUX_s_1_2_2(or_2742_cse, mux_tmp_824, fsm_output[5]);
  assign and_1055_ssc = and_dcpl_732 & and_dcpl_592;
  assign and_1059_ssc = and_dcpl_743 & and_dcpl_551 & and_dcpl_835;
  assign or_2741_nl = (~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1])
      | (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2) | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0])))
      | (~ (fsm_output[6])) | (fsm_output[8]);
  assign mux_2027_nl = MUX_s_1_2_2(or_tmp_464, mux_tmp_121, or_2739_cse);
  assign mux_2028_nl = MUX_s_1_2_2(or_2741_nl, mux_2027_nl, fsm_output[4]);
  assign mux_2029_nl = MUX_s_1_2_2(or_tmp_464, mux_2028_nl, fsm_output[0]);
  assign mux_2030_nl = MUX_s_1_2_2(mux_2029_nl, mux_tmp_824, fsm_output[5]);
  assign mux_2031_nl = MUX_s_1_2_2(mux_2030_nl, mux_2025_cse, fsm_output[1]);
  assign mux_2033_nl = MUX_s_1_2_2(mux_2032_cse, mux_2031_nl, and_1773_cse);
  assign APPLY_ROTARY_POS_EMB_LOOP_6_and_30_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (mux_2033_nl | (fsm_output[7]));
  assign and_1060_itm = and_dcpl_732 & and_dcpl_613;
  assign nor_410_nl = ~((~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd)
      | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1]) | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2
      | (~ (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0])));
  assign mux_2036_nl = MUX_s_1_2_2(mux_tmp_1945, mux_tmp_1943, nor_410_nl);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_and_18_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~((~ mux_2036_nl) & and_dcpl_259));
  assign and_1062_ssc = and_dcpl_732 & and_dcpl_607;
  assign and_1626_nl = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd & (~
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1])) & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2
      & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0]);
  assign mux_2037_nl = MUX_s_1_2_2(mux_tmp_1945, mux_tmp_1943, and_1626_nl);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_and_19_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~((~ mux_2037_nl) & and_dcpl_259));
  assign attention_2_1_16_16_4_4_k_proj_re_and_91_cse = (~ RESHAPE_2D_TO_3D_LOOP_2_2_and_cse)
      & and_dcpl_1034;
  assign attention_2_1_16_16_4_4_k_proj_re_or_cse = and_dcpl_1033 | attention_2_1_16_16_4_4_k_proj_re_and_91_cse;
  assign attention_2_1_16_16_4_4_k_proj_re_or_17_cse = (RESHAPE_2D_TO_3D_LOOP_2_2_and_cse
      & and_dcpl_1034) | and_dcpl_213;
  assign and_1771_cse = (fsm_output[2]) & (fsm_output[4]);
  assign mux_2087_nl = MUX_s_1_2_2(not_tmp_874, or_tmp_1132, fsm_output[7]);
  assign mux_2086_nl = MUX_s_1_2_2(not_tmp_874, or_tmp_1218, fsm_output[7]);
  assign mux_2088_nl = MUX_s_1_2_2(mux_2087_nl, mux_2086_nl, reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign nor_1228_ssc = ~(mux_2088_nl | (fsm_output[8]));
  assign nand_357_nl = ~((fsm_output[6]) & mux_tmp_1489);
  assign mux_1542_nl = MUX_s_1_2_2(nand_357_nl, or_tmp_1132, fsm_output[7]);
  assign attention_2_1_16_16_4_4_q_proj_and_5_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (mux_1542_nl | (fsm_output[8]) | and_dcpl_626);
  assign or_2792_cse = (fsm_output[1:0]!=2'b01);
  assign or_2797_cse = (fsm_output[4:3]!=2'b00);
  assign mux_2092_cse = MUX_s_1_2_2(or_2457_cse, or_1197_cse, fsm_output[4]);
  assign or_2799_nl = (~ (fsm_output[0])) | (fsm_output[1]) | (~ (fsm_output[4]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (fsm_output[8]);
  assign mux_2097_nl = MUX_s_1_2_2(or_2460_cse, or_tmp_1643, or_1732_cse);
  assign mux_2098_nl = MUX_s_1_2_2(or_2799_nl, mux_2097_nl, fsm_output[3]);
  assign mux_2096_nl = MUX_s_1_2_2(mux_1522_cse, or_1197_cse, or_2797_cse);
  assign mux_2099_nl = MUX_s_1_2_2(mux_2098_nl, mux_2096_nl, fsm_output[5]);
  assign mux_2093_nl = MUX_s_1_2_2(mux_2092_cse, or_tmp_1643, or_2792_cse);
  assign mux_2094_nl = MUX_s_1_2_2(or_2460_cse, mux_2093_nl, fsm_output[3]);
  assign or_2787_nl = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[4]);
  assign mux_2090_nl = MUX_s_1_2_2(mux_1522_cse, or_1197_cse, or_2787_nl);
  assign or_2786_nl = ((fsm_output[0]) & (fsm_output[1]) & (fsm_output[4])) | (fsm_output[8:6]!=3'b100);
  assign mux_2091_nl = MUX_s_1_2_2(mux_2090_nl, or_2786_nl, fsm_output[3]);
  assign mux_2095_nl = MUX_s_1_2_2(mux_2094_nl, mux_2091_nl, fsm_output[5]);
  assign mux_2100_ssc = MUX_s_1_2_2(mux_2099_nl, mux_2095_nl, fsm_output[2]);
  assign APPLY_ROTARY_POS_EMB_LOOP_6_and_28_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (and_dcpl_888 | and_dcpl_257 | and_dcpl_1073 | and_dcpl_240 | and_dcpl_207
      | and_dcpl_847 | and_dcpl_583);
  assign APPLY_ROTARY_POS_EMB_LOOP_6_and_31_cse = APPLY_ROTARY_POS_EMB_LOOP_6_and_28_cse
      & (~ and_dcpl_725);
  assign nand_283_nl = ~((fsm_output[6]) & mux_tmp_1421);
  assign mux_2102_nl = MUX_s_1_2_2(nand_283_nl, or_tmp_1218, fsm_output[7]);
  assign attention_2_1_16_16_4_4_q_proj_re_and_29_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (mux_2102_nl | (fsm_output[8]));
  assign mux_2103_nl = MUX_s_1_2_2((~ or_tmp_728), or_tmp_762, fsm_output[5]);
  assign mux_2104_nl = MUX_s_1_2_2(mux_tmp_91, mux_2103_nl, fsm_output[3]);
  assign attention_2_1_16_16_4_4_k_proj_re_and_65_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~((~ mux_2104_nl) & and_dcpl_259));
  assign attention_2_1_16_16_4_4_v_proj_re_and_32_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~(((and_1638_cse | (fsm_output[4])) ^ (fsm_output[5])) & and_dcpl_259));
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_and_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~((~ (fsm_output[2])) | (fsm_output[4]) | (fsm_output[8]) | nand_197_cse
      | or_dcpl_1134 | or_1983_cse));
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_and_29_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (and_dcpl_257 | and_dcpl_410 | and_dcpl_240 | and_dcpl_1034 | and_dcpl_207
      | and_dcpl_213 | and_dcpl_583 | and_dcpl_265);
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse = and_dcpl_410 | attention_2_1_16_16_4_4_k_proj_re_and_91_cse;
  assign nand_285_nl = ~((fsm_output[6]) & mux_tmp_857);
  assign or_2828_nl = (fsm_output[5]) | nor_tmp_282;
  assign mux_2107_nl = MUX_s_1_2_2(or_2828_nl, or_2699_cse, fsm_output[3]);
  assign or_3153_nl = (fsm_output[6]) | mux_2107_nl;
  assign mux_2108_nl = MUX_s_1_2_2(nand_285_nl, or_3153_nl, fsm_output[7]);
  assign attention_2_1_16_16_4_4_v_proj_re_and_95_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (mux_2108_nl | (fsm_output[8]));
  assign mux_2109_nl = MUX_s_1_2_2(nor_717_cse, or_3137_cse, fsm_output[3]);
  assign attention_2_1_16_16_4_4_v_proj_and_30_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~((~(mux_2109_nl | (fsm_output[8]))) & and_dcpl_1145));
  assign GEMM_3D_FLOAT_LOOP_3_1_mux_4_nl = MUX_s_1_2_2((~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1),
      (~ or_dcpl_1155), and_dcpl_1154);
  assign mux_2124_nl = MUX_s_1_2_2(nand_tmp_99, or_tmp_1664, or_270_cse);
  assign mux_2123_nl = MUX_s_1_2_2(mux_tmp_2116, or_tmp_1671, fsm_output[2]);
  assign mux_2125_nl = MUX_s_1_2_2(mux_2124_nl, mux_2123_nl, fsm_output[3]);
  assign mux_2126_nl = MUX_s_1_2_2(mux_2125_nl, mux_tmp_2121, fsm_output[1]);
  assign or_2840_nl = (fsm_output[8:5]!=4'b1000);
  assign mux_2114_nl = MUX_s_1_2_2(or_tmp_1664, or_2840_nl, and_1771_cse);
  assign mux_2120_nl = MUX_s_1_2_2(mux_tmp_2119, mux_2114_nl, fsm_output[3]);
  assign mux_2122_nl = MUX_s_1_2_2(mux_tmp_2121, mux_2120_nl, fsm_output[1]);
  assign mux_2127_nl = MUX_s_1_2_2(mux_2126_nl, mux_2122_nl, fsm_output[0]);
  assign GEMM_3D_FLOAT_LOOP_3_1_and_44_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((GEMM_3D_FLOAT_LOOP_3_1_mux_4_nl & mux_2127_nl) | and_dcpl_1152 | and_dcpl_222);
  assign mux_2128_nl = MUX_s_1_2_2(or_3167_cse, or_1907_cse, fsm_output[0]);
  assign attention_2_1_16_16_4_4_q_embed_and_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~((~ mux_2128_nl) & and_dcpl_201 & and_dcpl_199));
  assign and_1782_cse = (fsm_output[4:2]==3'b111);
  assign nor_1239_cse = ~((fsm_output[5]) | and_1782_cse | (fsm_output[6]) | (~ (fsm_output[8])));
  assign nor_593_cse = ~((fsm_output[2:1]!=2'b01));
  assign nor_1240_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_1241_nl = ~((~((fsm_output[4]) | (fsm_output[6]))) | (fsm_output[8]));
  assign mux_2155_nl = MUX_s_1_2_2(nor_1240_nl, nor_1241_nl, and_1474_cse);
  assign nor_1242_nl = ~((~((~((fsm_output[1]) | (fsm_output[0]) | (~ (fsm_output[4]))))
      | (fsm_output[6]))) | (fsm_output[8]));
  assign mux_2156_nl = MUX_s_1_2_2(mux_2155_nl, nor_1242_nl, fsm_output[2]);
  assign nor_1243_nl = ~((~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_1244_nl = ~((~((~((fsm_output[0]) | (z_out_5[2]))) | (fsm_output[4])))
      | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_2154_nl = MUX_s_1_2_2(nor_1243_nl, nor_1244_nl, nor_593_cse);
  assign mux_2157_cse = MUX_s_1_2_2(mux_2156_nl, mux_2154_nl, fsm_output[3]);
  assign attention_2_1_16_16_4_4_attn_weights_and_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~(and_dcpl_185 & or_1732_cse & and_dcpl_190));
  assign GEMM_3D_FLOAT_LOOP_3_and_36_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~((or_1732_cse ^ (fsm_output[2])) & and_dcpl_61 & and_dcpl_190));
  assign attention_2_1_16_16_4_4_attn_weights_and_52_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~(and_dcpl_61 & (~ (fsm_output[2])) & (fsm_output[5]) & and_dcpl_1141));
  assign attention_2_1_16_16_4_4_attn_weights_and_48_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~ and_dcpl_1195);
  assign mux_1543_nl = MUX_s_1_2_2((~ (fsm_output[2])), (fsm_output[2]), fsm_output[1]);
  assign mux_2237_nl = MUX_s_1_2_2(or_3167_cse, mux_1543_nl, fsm_output[0]);
  assign attention_2_1_16_16_4_4_attn_weights_and_12_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~((~ mux_2237_nl) & and_dcpl_61 & and_dcpl_293));
  assign attention_2_1_16_16_4_4_attn_weights_and_24_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~ and_dcpl_304);
  assign GEMM_3D_FLOAT_LOOP_3_1_and_46_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~((~(mux_tmp_1440 | (fsm_output[8]))) & nor_646_cse & and_dcpl_148));
  assign mux_2249_nl = MUX_s_1_2_2((~ nor_tmp_285), or_tmp_861, fsm_output[5]);
  assign mux_2250_nl = MUX_s_1_2_2(mux_2249_nl, or_tmp_682, fsm_output[3]);
  assign attention_abs_4_qelse_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~((~ mux_2250_nl) & and_dcpl_258 & (fsm_output[7])));
  assign compute_sqrt_1_guess_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((and_dcpl_362 & and_dcpl_221) | and_dcpl_292);
  assign attention_2_1_16_16_4_4_quantized_final_output_and_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1158 | (~ mux_2256_itm))) | mux_tmp_2252);
  assign RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse = (~ QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1)
      & and_dcpl_1154;
  assign RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse = QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1
      & and_dcpl_1154;
  assign attention_2_1_16_16_4_4_quantized_final_output_and_8_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1166 | (~ mux_2256_itm))) | mux_tmp_2252);
  assign attention_2_1_16_16_4_4_quantized_final_output_and_16_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1164 | (~ mux_2256_itm))) | mux_tmp_2252);
  assign attention_2_1_16_16_4_4_quantized_final_output_and_24_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1161 | (~ mux_2256_itm))) | mux_tmp_2252);
  assign attention_2_1_16_16_4_4_quantized_final_output_and_32_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1159 | (~ mux_2256_itm))) | mux_tmp_2252);
  assign attention_2_1_16_16_4_4_quantized_final_output_and_40_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1156 | (~ mux_2256_itm))) | mux_tmp_2252);
  assign attention_2_1_16_16_4_4_quantized_final_output_and_48_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1160 | (~ mux_2256_itm))) | mux_tmp_2252);
  assign attention_2_1_16_16_4_4_quantized_final_output_and_56_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1162 | (~ mux_2256_itm))) | mux_tmp_2252);
  assign attention_2_1_16_16_4_4_quantized_final_output_and_64_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1165 | (~ mux_2256_itm))) | mux_tmp_2252);
  assign attention_2_1_16_16_4_4_quantized_final_output_and_72_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1167 | (~ mux_2256_itm))) | mux_tmp_2252);
  assign attention_2_1_16_16_4_4_quantized_final_output_and_80_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1169 | (~ mux_2256_itm))) | mux_tmp_2252);
  assign attention_2_1_16_16_4_4_quantized_final_output_and_88_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1141 | (~ mux_2256_itm))) | mux_tmp_2252);
  assign attention_2_1_16_16_4_4_quantized_final_output_and_96_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1170 | (~ mux_2256_itm))) | mux_tmp_2252);
  assign attention_2_1_16_16_4_4_quantized_final_output_and_104_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & ((~(or_dcpl_1168 | (~ mux_2256_itm))) | mux_tmp_2252);
  assign mux_2257_nl = MUX_s_1_2_2(or_dcpl_1050, nor_tmp_329, fsm_output[5]);
  assign mux_2258_nl = MUX_s_1_2_2((fsm_output[5]), (~ mux_2257_nl), fsm_output[3]);
  assign attention_2_1_16_16_4_4_quantized_final_output_and_112_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (~(mux_2258_nl & and_dcpl_413));
  assign attention_2_1_16_16_4_4_v_proj_re_and_63_cse = (~ or_dcpl_1141) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_65_cse = (~ or_dcpl_1170) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_67_cse = (~ or_dcpl_1169) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_69_cse = (~ or_dcpl_1168) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_71_cse = (~ or_dcpl_1167) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_73_cse = (~ or_dcpl_1166) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_75_cse = (~ or_dcpl_1165) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_77_cse = (~ or_dcpl_1164) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_79_cse = (~ or_dcpl_1162) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_81_cse = (~ or_dcpl_1161) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_83_cse = (~ or_dcpl_1160) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_85_cse = (~ or_dcpl_1159) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_87_cse = (~ or_dcpl_1158) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_89_cse = (~ or_dcpl_1156) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_91_cse = (~ or_dcpl_1155) & and_dcpl_1225;
  assign attention_2_1_16_16_4_4_v_proj_re_and_93_cse = (~ or_dcpl_1152) & and_dcpl_1225;
  assign output_and_16_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 &
      (~(((and_1771_cse & (fsm_output[1]) & (fsm_output[3])) ^ (fsm_output[5])) &
      and_dcpl_413));
  assign output_and_64_cse = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 &
      (~ and_dcpl_1232);
  assign or_1659_nl = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd | (~ GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva);
  assign attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2_mx1 = MUX_v_40_2_2(acc_3_cse_40_1,
      attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3, or_1659_nl);
  assign nand_298_nl = ~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0);
  assign attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2_mx1 = MUX_v_40_2_2(acc_3_cse_40_1,
      attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3, nand_298_nl);
  assign or_1661_nl = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd | (~ GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva);
  assign attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2_mx1 = MUX_v_40_2_2(acc_3_cse_40_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2, or_1661_nl);
  assign nand_299_nl = ~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  assign attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2_mx1 = MUX_v_40_2_2(acc_3_cse_40_1,
      attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3, nand_299_nl);
  assign or_1663_nl = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd | (~ GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva);
  assign attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2_mx1 = MUX_v_40_2_2(acc_3_cse_40_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2, or_1663_nl);
  assign nand_300_nl = ~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva);
  assign attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2_mx1 = MUX_v_40_2_2(acc_3_cse_40_1,
      attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3, nand_300_nl);
  assign or_1665_nl = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd | (~ GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva);
  assign attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2_mx1 = MUX_v_40_2_2(acc_3_cse_40_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2, or_1665_nl);
  assign nand_301_nl = ~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd & GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva);
  assign attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2_mx1 = MUX_v_40_2_2(acc_3_cse_40_1,
      attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3, nand_301_nl);
  assign or_1667_ssc = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd | (~ GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva);
  assign attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_39 = MUX_s_1_2_2((acc_3_cse_40_1[39]),
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd, or_1667_ssc);
  assign attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_38_0 = MUX_v_39_2_2((acc_3_cse_40_1[38:0]),
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1, or_1667_ssc);
  assign or_1669_nl = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd | (~ GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva);
  assign attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2_mx1 = MUX_v_40_2_2(acc_3_cse_40_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2, or_1669_nl);
  assign or_1671_nl = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd | (~ reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  assign attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2_mx1 = MUX_v_40_2_2(acc_3_cse_40_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2, or_1671_nl);
  assign attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2_mx1 = MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva);
  assign attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2_mx1 = MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_1,
      acc_3_cse_40_1, reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  assign attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2_mx1 = MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva);
  assign attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2_mx1 = MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_1,
      acc_3_cse_40_1, LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0);
  assign attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2_mx1 = MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva);
  assign attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2_mx1 = MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva);
  assign attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2_mx1 = MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva);
  assign attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2_mx1 = MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva);
  assign attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2_mx1 = MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva);
  assign attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2_mx1 = MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva);
  assign attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2_mx1 = MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva);
  assign attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2_mx1 = MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_1,
      acc_3_cse_40_1, GEMM_3D_FLOAT_LOOP_3_and_tmp_sva);
  assign attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1, or_dcpl_980);
  assign attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1, or_dcpl_983);
  assign attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1, or_dcpl_985);
  assign attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1, or_dcpl_989);
  assign attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1, or_dcpl_990);
  assign attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1, or_dcpl_993);
  assign attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1, or_dcpl_998);
  assign attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3, or_dcpl_980);
  assign attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3, or_dcpl_983);
  assign attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3, or_dcpl_985);
  assign attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3, or_dcpl_987);
  assign attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2, or_dcpl_988);
  assign attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3, or_dcpl_989);
  assign and_1455_cse = (((fsm_output[4]) & (fsm_output[6])) | (fsm_output[7])) &
      (fsm_output[8]);
  assign nor_176_cse = ~((fsm_output[1]) | (~ (fsm_output[4])));
  assign attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2, or_dcpl_990);
  assign attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2, or_dcpl_993);
  assign attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2, or_dcpl_996);
  assign attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2, or_dcpl_998);
  assign attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1, or_dcpl_1000);
  assign attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_39_16, or_dcpl_1002);
  assign attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0_mx0w1 = MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_15_0, or_dcpl_1002);
  assign attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_39_16, or_dcpl_1004);
  assign attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0_mx0w1 = MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_15_0, or_dcpl_1004);
  assign attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_39_16, or_dcpl_1006);
  assign attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0_mx0w1 = MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_15_0, or_dcpl_1006);
  assign attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16, or_dcpl_1008);
  assign attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0_mx0w1 = MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_15_0, or_dcpl_1008);
  assign attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_39_16, or_dcpl_1009);
  assign attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0_mx0w1 = MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_15_0, or_dcpl_1009);
  assign attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16, or_dcpl_1010);
  assign attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_39_16, or_dcpl_1011);
  assign attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0_mx0w1 = MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_15_0, or_dcpl_1011);
  assign attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16, or_dcpl_1012);
  assign attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_39_16, or_dcpl_1013);
  assign attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0_mx0w1 = MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0, or_dcpl_1013);
  assign attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16, or_dcpl_1014);
  assign attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_39_16, or_dcpl_1015);
  assign attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0_mx0w1 = MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_15_0, or_dcpl_1015);
  assign attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16, or_dcpl_1016);
  assign attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_39_16, or_dcpl_1017);
  assign attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0_mx0w1 = MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_15_0, or_dcpl_1017);
  assign attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16, or_dcpl_1018);
  assign attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16, or_dcpl_1019);
  assign attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0_mx0w1 = MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_15_0, or_dcpl_1019);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2, or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2, or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w0 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2, or_dcpl_1023);
  assign mux_502_cse = MUX_s_1_2_2(or_2456_cse, (fsm_output[8]), fsm_output[7]);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w3 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2, or_dcpl_1025);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2_mx0w1 = MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16_mx0w1 = MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1,
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 =
      MUX_v_8_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm,
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm,
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16_mx0w1 = MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_39_16, or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_13
      = MUX_v_3_2_2((APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm[7:5]),
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd, or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_12_8 =
      MUX_v_5_2_2((APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm[4:0]),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1[12:8]),
      or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1[7]), or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1[6]), or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1[5]), or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1[4]), or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1[3]), or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1[2]), or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1[1]), or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm,
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1[0]), or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16_mx0w1 = MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_39_16, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 =
      MUX_v_8_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_15_8, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_7, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_6, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_5, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_4, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_3, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_2, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_1, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_0, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 =
      MUX_v_8_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0, or_dcpl_1023);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16_mx0w1 = MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16, or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 =
      MUX_v_8_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd, or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7, or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6, or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5, or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4, or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3, or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2, or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1, or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0, or_dcpl_1021);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16_mx0w1 = MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_39_16, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8 =
      MUX_v_8_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1, or_dcpl_1024);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0 = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0, or_dcpl_1024);
  assign attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out[15:8]),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_15_8, or_dcpl_1028);
  assign attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out[7]),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7, or_dcpl_1028);
  assign attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out[6]),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6, or_dcpl_1028);
  assign attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out[5]),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5, or_dcpl_1028);
  assign attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out[4]),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4, or_dcpl_1028);
  assign attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out[3]),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3, or_dcpl_1028);
  assign attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out[2]),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2, or_dcpl_1028);
  assign attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out[1]),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1, or_dcpl_1028);
  assign attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out[0]),
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0, or_dcpl_1028);
  assign attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out[15:8]),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_15_8, or_dcpl_1030);
  assign attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out[7]),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7, or_dcpl_1030);
  assign attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out[6]),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6, or_dcpl_1030);
  assign attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out[5]),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5, or_dcpl_1030);
  assign attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out[4]),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4, or_dcpl_1030);
  assign attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out[3]),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3, or_dcpl_1030);
  assign attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out[2]),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2, or_dcpl_1030);
  assign attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out[1]),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1, or_dcpl_1030);
  assign attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out[0]),
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0, or_dcpl_1030);
  assign attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out[15:8]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_15_8, or_dcpl_1031);
  assign attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out[7]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7, or_dcpl_1031);
  assign attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out[6]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6, or_dcpl_1031);
  assign attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out[5]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5, or_dcpl_1031);
  assign attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out[4]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4, or_dcpl_1031);
  assign attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out[3]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3, or_dcpl_1031);
  assign attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out[2]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2, or_dcpl_1031);
  assign attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out[1]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1, or_dcpl_1031);
  assign attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out[0]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0, or_dcpl_1031);
  assign attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out[15:8]),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_15_8, or_dcpl_1033);
  assign attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out[7]),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7, or_dcpl_1033);
  assign attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out[6]),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6, or_dcpl_1033);
  assign attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out[5]),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5, or_dcpl_1033);
  assign attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out[4]),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4, or_dcpl_1033);
  assign attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out[3]),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3, or_dcpl_1033);
  assign attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out[2]),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2, or_dcpl_1033);
  assign attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out[1]),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1, or_dcpl_1033);
  assign attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out[0]),
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0, or_dcpl_1033);
  assign attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out[15:8]),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_15_8, or_dcpl_1035);
  assign attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out[7]),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7, or_dcpl_1035);
  assign attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out[6]),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6, or_dcpl_1035);
  assign attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out[5]),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5, or_dcpl_1035);
  assign attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out[4]),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4, or_dcpl_1035);
  assign attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out[3]),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3, or_dcpl_1035);
  assign attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out[2]),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2, or_dcpl_1035);
  assign attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out[1]),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1, or_dcpl_1035);
  assign attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out[0]),
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0, or_dcpl_1035);
  assign attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out[15:8]),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_15_8, or_dcpl_1037);
  assign attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out[7]),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7, or_dcpl_1037);
  assign attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out[6]),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6, or_dcpl_1037);
  assign attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out[5]),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5, or_dcpl_1037);
  assign attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out[4]),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4, or_dcpl_1037);
  assign attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out[3]),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3, or_dcpl_1037);
  assign attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out[2]),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2, or_dcpl_1037);
  assign attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out[1]),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1, or_dcpl_1037);
  assign attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out[0]),
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0, or_dcpl_1037);
  assign attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out[15:8]),
      attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_8, or_dcpl_1038);
  assign attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out[7]),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd, or_dcpl_1038);
  assign attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out[6]),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_1, or_dcpl_1038);
  assign attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out[5]),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_2, or_dcpl_1038);
  assign attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out[4]),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_3, or_dcpl_1038);
  assign attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out[3]),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_4, or_dcpl_1038);
  assign attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out[2]),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_5, or_dcpl_1038);
  assign attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out[1]),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_6, or_dcpl_1038);
  assign attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out[0]),
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_7, or_dcpl_1038);
  assign attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out[15:8]),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_15_8, or_dcpl_1039);
  assign attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out[7]),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_7, or_dcpl_1039);
  assign attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out[6]),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_6, or_dcpl_1039);
  assign attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out[5]),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_5, or_dcpl_1039);
  assign attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out[4]),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_4, or_dcpl_1039);
  assign attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out[3]),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_3, or_dcpl_1039);
  assign attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out[2]),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_2, or_dcpl_1039);
  assign attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out[1]),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_1, or_dcpl_1039);
  assign attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out[0]),
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_0, or_dcpl_1039);
  assign attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out[15:8]),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_15_8, or_dcpl_1041);
  assign attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out[7]),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7, or_dcpl_1041);
  assign attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out[6]),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6, or_dcpl_1041);
  assign attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out[5]),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5, or_dcpl_1041);
  assign attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out[4]),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4, or_dcpl_1041);
  assign attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out[3]),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3, or_dcpl_1041);
  assign attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out[2]),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2, or_dcpl_1041);
  assign attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out[1]),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1, or_dcpl_1041);
  assign attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out[0]),
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0, or_dcpl_1041);
  assign attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0_mx0w1 = MUX_v_16_2_2(z_out,
      attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_15_0, or_dcpl_1042);
  assign attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out[15:8]),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_15_8, or_dcpl_1043);
  assign attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out[7]),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7, or_dcpl_1043);
  assign attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out[6]),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6, or_dcpl_1043);
  assign attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out[5]),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5, or_dcpl_1043);
  assign attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out[4]),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4, or_dcpl_1043);
  assign attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out[3]),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3, or_dcpl_1043);
  assign attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out[2]),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2, or_dcpl_1043);
  assign attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out[1]),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1, or_dcpl_1043);
  assign attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out[0]),
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0, or_dcpl_1043);
  assign attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0_mx0w1 = MUX_v_16_2_2(z_out,
      attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_15_0, or_dcpl_1044);
  assign attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out[15:8]),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_15_8, or_dcpl_1045);
  assign attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out[7]),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7, or_dcpl_1045);
  assign attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out[6]),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6, or_dcpl_1045);
  assign attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out[5]),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5, or_dcpl_1045);
  assign attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out[4]),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4, or_dcpl_1045);
  assign attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out[3]),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3, or_dcpl_1045);
  assign attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out[2]),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2, or_dcpl_1045);
  assign attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out[1]),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1, or_dcpl_1045);
  assign attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out[0]),
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0, or_dcpl_1045);
  assign attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out[15:8]),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_15_8, or_dcpl_1046);
  assign attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out[7]),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7, or_dcpl_1046);
  assign attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out[6]),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6, or_dcpl_1046);
  assign attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out[5]),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5, or_dcpl_1046);
  assign attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out[4]),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4, or_dcpl_1046);
  assign attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out[3]),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3, or_dcpl_1046);
  assign attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out[2]),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2, or_dcpl_1046);
  assign attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out[1]),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1, or_dcpl_1046);
  assign attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out[0]),
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0, or_dcpl_1046);
  assign attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16, or_dcpl_1002);
  assign attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out_1[15:8]),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_15_8, or_dcpl_1002);
  assign attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out_1[7]),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_7, or_dcpl_1002);
  assign attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out_1[6]),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_6, or_dcpl_1002);
  assign attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out_1[5]),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_5, or_dcpl_1002);
  assign attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out_1[4]),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_4, or_dcpl_1002);
  assign attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out_1[3]),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_3, or_dcpl_1002);
  assign attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out_1[2]),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_2, or_dcpl_1002);
  assign attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out_1[1]),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_1, or_dcpl_1002);
  assign attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out_1[0]),
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_0, or_dcpl_1002);
  assign attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_39_16, or_dcpl_1004);
  assign attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0_mx0w1 = MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0, or_dcpl_1004);
  assign attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_39_16, or_dcpl_1006);
  assign attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_15_13 = MUX_v_3_2_2((z_out_1[15:13]),
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd, or_dcpl_1006);
  assign attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0 = MUX_v_13_2_2((z_out_1[12:0]),
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1, or_dcpl_1006);
  assign attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_39_16, or_dcpl_1008);
  assign attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0_mx0w1 = MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_15_0, or_dcpl_1008);
  assign attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_39_16, or_dcpl_1009);
  assign attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0_mx0w1 = MUX_v_16_2_2(z_out_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0, or_dcpl_1009);
  assign attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_39_16, or_dcpl_1010);
  assign attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0_mx0w1 = MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_15_0, or_dcpl_1010);
  assign attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48, or_dcpl_1011);
  assign attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_39_16, or_dcpl_1012);
  assign attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0_mx0w1 = MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0, or_dcpl_1012);
  assign attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_39_16, or_dcpl_1013);
  assign attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out_1[15:8]),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8, or_dcpl_1013);
  assign attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out_1[7]),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7, or_dcpl_1013);
  assign attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out_1[6]),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6, or_dcpl_1013);
  assign attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out_1[5]),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5, or_dcpl_1013);
  assign attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out_1[4]),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4, or_dcpl_1013);
  assign attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out_1[3]),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3, or_dcpl_1013);
  assign attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out_1[2]),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2, or_dcpl_1013);
  assign attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out_1[1]),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1, or_dcpl_1013);
  assign attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out_1[0]),
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0, or_dcpl_1013);
  assign attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_39_16, or_dcpl_1014);
  assign attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0_mx0w1 = MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_15_0, or_dcpl_1014);
  assign attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16, or_dcpl_1015);
  assign attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out_1[15:8]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd, or_dcpl_1015);
  assign attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out_1[7]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7, or_dcpl_1015);
  assign attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out_1[6]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6, or_dcpl_1015);
  assign attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out_1[5]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5, or_dcpl_1015);
  assign attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out_1[4]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4, or_dcpl_1015);
  assign attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out_1[3]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3, or_dcpl_1015);
  assign attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out_1[2]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2, or_dcpl_1015);
  assign attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out_1[1]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1, or_dcpl_1015);
  assign attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out_1[0]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0, or_dcpl_1015);
  assign attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_39_16, or_dcpl_1016);
  assign attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0_mx0w1 = MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_15_0, or_dcpl_1016);
  assign attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_15_8 = MUX_v_8_2_2((z_out_1[15:8]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd, or_dcpl_1017);
  assign attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_7 = MUX_s_1_2_2((z_out_1[7]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7, or_dcpl_1017);
  assign attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_6 = MUX_s_1_2_2((z_out_1[6]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6, or_dcpl_1017);
  assign attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_5 = MUX_s_1_2_2((z_out_1[5]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5, or_dcpl_1017);
  assign attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_4 = MUX_s_1_2_2((z_out_1[4]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4, or_dcpl_1017);
  assign attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_3 = MUX_s_1_2_2((z_out_1[3]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3, or_dcpl_1017);
  assign attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_2 = MUX_s_1_2_2((z_out_1[2]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2, or_dcpl_1017);
  assign attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_1 = MUX_s_1_2_2((z_out_1[1]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1, or_dcpl_1017);
  assign attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_0 = MUX_s_1_2_2((z_out_1[0]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0, or_dcpl_1017);
  assign attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_39_16, or_dcpl_1018);
  assign attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0_mx0w1 = MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_15_0, or_dcpl_1018);
  assign attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16_mx0w1 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_39_16, or_dcpl_1019);
  assign attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0_mx0w1 = MUX_v_16_2_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_15_0, or_dcpl_1019);
  assign nor_749_cse = ~((fsm_output[2]) | (fsm_output[0]));
  assign or_76_cse = reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 | reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd;
  assign or_130_cse = (~ reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1) | reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd;
  assign drf_output_sdt_2_sva_15_0_mx0w0 = MUX_v_16_16_2(attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0,
      ({APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8 , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6 , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4 , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2 , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0}), attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_15_0,
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0, attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_15_0,
      attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_15_0, attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_15_0,
      attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0, attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_15_0,
      attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_15_0, ({reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd
      , reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1}), ({apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_15_8
      , apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_7 , apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_6
      , apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_5 , apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_4
      , apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_3 , apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_2
      , apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_1 , apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_0}),
      attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0, attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_15_0,
      attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_15_0, attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0,
      {reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2});
  assign drf_output_sdt_3_sva_15_0_mx0w3 = MUX_v_16_16_2(attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0,
      ({APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8 , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6 , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4 , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2 , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0}), apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0,
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0, attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0, {reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2});
  assign SOFTMAX_LOOP_5_mux_12_psp_mx0w0 = MUX_v_40_12_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_5,
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_5, attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_5,
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_5, attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_4,
      attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_4, attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_4,
      attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_4, attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_4,
      attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_4, attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_4,
      attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_4, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_2_conc_1_mut_71_48_mx0w0 = MUX_v_24_16_2(attention_2_1_16_16_4_4_v_proj_re_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_3_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_4_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_5_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_6_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_7_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_8_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_9_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_10_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_12_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_13_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_14_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_15_sva_1_39_16, {reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2});
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_3_conc_1_mut_71_48_mx0w3 = MUX_v_24_16_2(output_0_0_sva_1_39_16,
      output_0_1_sva_1_39_16, output_0_2_sva_1_39_16, output_0_3_sva_1_39_16, output_0_4_sva_1_39_16,
      output_0_5_sva_1_39_16, output_0_6_sva_1_39_16, output_0_7_sva_1_39_16, output_0_8_sva_1_39_16,
      output_0_9_sva_1_39_16, output_0_10_sva_1_39_16, output_0_11_sva_1_39_16, output_0_12_sva_1_39_16,
      output_0_13_sva_1_39_16, output_0_14_sva_1_39_16, output_0_15_sva_1_39_16,
      {reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2});
  assign nl_compute_sqrt_1_for_acc_1_nl = conv_s2s_40_41({LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4
      , LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0 , compute_sqrt_1_guess_sva_34
      , compute_sqrt_1_guess_sva_33_0}) + conv_s2s_40_41(APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm[39:0]);
  assign compute_sqrt_1_for_acc_1_nl = nl_compute_sqrt_1_for_acc_1_nl[40:0];
  assign compute_sqrt_1_for_acc_1_itm_40_1_1 = readslicef_41_40_1(compute_sqrt_1_for_acc_1_nl);
  assign nl_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2 = $signed(GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm)
      * $signed(22'b0100101101010110010011);
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2 = nl_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2[60:0];
  assign or_1860_nl = reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 | (CM_LOOP_3_acc_tmp[0]);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx1 = MUX_v_40_2_2(CM_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_ctmp_sva_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_3, or_1860_nl);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx2 = MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z[39:0]),
      attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_5, or_dcpl_1063);
  assign attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_39 =
      reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 & attention_max_attn_fixed_t_1_acc_1_itm_40_1;
  assign attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_38_0
      = MUX_v_39_2_2(39'b000000000000000000000000000000000000000, reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1,
      attention_max_attn_fixed_t_1_acc_1_itm_40_1);
  assign nl_compute_sqrt_for_acc_1_nl = conv_s2s_40_41({LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4
      , LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0 , compute_sqrt_guess_sva_34
      , compute_sqrt_guess_sva_33_0}) + conv_s2s_40_41(APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm[39:0]);
  assign compute_sqrt_for_acc_1_nl = nl_compute_sqrt_for_acc_1_nl[40:0];
  assign compute_sqrt_for_acc_1_itm_40_1_1 = readslicef_41_40_1(compute_sqrt_for_acc_1_nl);
  assign nl_attention_abs_1_qr_sva_1 = conv_u2s_39_40(~ (input_0_0_sva_2[38:0]))
      + 40'b0000000000000000000000000000000000000001;
  assign attention_abs_1_qr_sva_1 = nl_attention_abs_1_qr_sva_1[39:0];
  assign nl_softmax_1_4_3_sum_sva_2 = ({reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd , reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1})
      + SOFTMAX_LOOP_4_acc_3_cse_sva_1;
  assign softmax_1_4_3_sum_sva_2 = nl_softmax_1_4_3_sum_sva_2[39:0];
  assign attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx2 = MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z[39:0]),
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_5, or_dcpl_1076);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx1 = MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z[39:0]),
      attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_4, or_dcpl_1081);
  assign nl_LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp = conv_u2s_4_5({reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2})
      + 5'b00001;
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp = nl_LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp[4:0];
  assign nl_RMS_NORM_LOOP_2_2_acc_1_tmp = conv_u2s_4_5({reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
      , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1}) + 5'b00001;
  assign RMS_NORM_LOOP_2_2_acc_1_tmp = nl_RMS_NORM_LOOP_2_2_acc_1_tmp[4:0];
  assign nl_attention_abs_qr_35_0_lpi_1_dfm_mx0w0 = conv_u2s_35_36(~ (operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1[34:0]))
      + 36'b000000000000000000000000000000000001;
  assign attention_abs_qr_35_0_lpi_1_dfm_mx0w0 = nl_attention_abs_qr_35_0_lpi_1_dfm_mx0w0[35:0];
  assign attention_abs_qr_35_0_lpi_1_dfm_mx1_35 = (attention_abs_qr_35_0_lpi_1_dfm_mx0w0[35])
      & (operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1[35]);
  assign attention_abs_qr_35_0_lpi_1_dfm_mx1_34_1 = MUX_v_34_2_2((operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1[34:1]),
      (attention_abs_qr_35_0_lpi_1_dfm_mx0w0[34:1]), operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1[35]);
  assign operator_40_24_true_AC_TRN_AC_WRAP_and_1_nl = reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd
      & reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  assign nl_operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1
      = ({reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd , (reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[38:4])})
      + conv_u2s_1_36(operator_40_24_true_AC_TRN_AC_WRAP_and_1_nl);
  assign operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1
      = nl_operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1[35:0];
  assign QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_dfm_1_38_0_1 = MUX1HOT_v_39_5_2((input_0_0_sva_2[38:0]),
      reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1, QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_38_0,
      (RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva[38:0]), attention_abs_3_qr_sva_38_0,
      {RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_nor_1_ssc_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , RMS_NORM_LOOP_2_and_29_ssc , RMS_NORM_LOOP_2_and_33_ssc_1 , RMS_NORM_LOOP_2_and_34_ssc});
  assign RMS_NORM_LOOP_2_2_unequal_tmp_mx0w0 = ~(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4
      & (LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0==4'b1111));
  assign nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3 = conv_u2u_2_3(z_out_11[2:1])
      + conv_u2u_2_3({reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3 = nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3[2:0];
  assign nl_GEMM_3D_FLOAT_LOOP_3_acc_6_tmp = conv_u2u_2_3(z_out_11[2:1]) + conv_u2u_2_3({reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign GEMM_3D_FLOAT_LOOP_3_acc_6_tmp = nl_GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2:0];
  assign nl_attention_abs_2_mux_2 = conv_u2s_39_40(~ (RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva[38:0]))
      + 40'b0000000000000000000000000000000000000001;
  assign attention_abs_2_mux_2 = nl_attention_abs_2_mux_2[39:0];
  assign QUANTIZE_ACTIVATION_LOOP_2_attention_abs_2_nand_nl = ~((attention_abs_2_mux_2[39])
      & (RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva[39]));
  assign attention_abs_2_mux_3_nl = MUX_v_39_2_2((RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva[38:0]),
      (attention_abs_2_mux_2[38:0]), RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva[39]);
  assign nl_QUANTIZE_ACTIVATION_LOOP_2_acc_4_nl = conv_s2u_40_41({reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      , QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_38_0}) + conv_s2u_40_41({QUANTIZE_ACTIVATION_LOOP_2_attention_abs_2_nand_nl
      , (~ attention_abs_2_mux_3_nl)}) + 41'b00000000000000000000000000000000000000001;
  assign QUANTIZE_ACTIVATION_LOOP_2_acc_4_nl = nl_QUANTIZE_ACTIVATION_LOOP_2_acc_4_nl[40:0];
  assign QUANTIZE_ACTIVATION_LOOP_2_acc_4_itm_40_1 = readslicef_41_1_40(QUANTIZE_ACTIVATION_LOOP_2_acc_4_nl);
  assign RMS_NORM_LOOP_2_and_29_ssc_1 = (~ QUANTIZE_ACTIVATION_LOOP_2_acc_4_itm_40_1)
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign RMS_NORM_LOOP_2_and_34_ssc_1 = (RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva[39])
      & RMS_NORM_LOOP_2_and_30_m1c_1;
  assign RMS_NORM_LOOP_2_and_30_m1c_1 = QUANTIZE_ACTIVATION_LOOP_2_acc_4_itm_40_1
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign RMS_NORM_LOOP_2_2_and_32_ssc_mx0w3 = (attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_2_mx0[39])
      & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_nor_1_ssc_1 = ~((input_0_0_sva_2[39]) |
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign RMS_NORM_LOOP_2_and_33_ssc_1 = (~ (RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva[39]))
      & RMS_NORM_LOOP_2_and_30_m1c;
  assign QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_dfm_1_38_0_mx0w1 = MUX1HOT_v_39_5_2((attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1[38:0]),
      attention_abs_5_qr_sva_38_0, QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_38_0,
      (RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva[38:0]), attention_abs_7_qr_sva_38_0,
      {RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_nor_1_ssc_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , RMS_NORM_LOOP_2_2_and_29_ssc , RMS_NORM_LOOP_2_2_and_33_ssc_1 , RMS_NORM_LOOP_2_2_and_34_ssc});
  assign QUANTIZE_ACTIVATION_LOOP_3_nand_seb = ~((reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1==2'b11)
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd);
  assign QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse
      = ~(QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1 | QUANTIZE_ACTIVATION_LOOP_3_nand_seb);
  assign attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16, or_dcpl_1137);
  assign attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16, or_dcpl_1138);
  assign attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16, or_dcpl_1084);
  assign attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16, or_dcpl_1092);
  assign attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16, or_dcpl_1079);
  assign attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16, or_dcpl_1141);
  assign nl_QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_nl = ({1'b1 ,
      reg_QUANTIZE_ACTIVATION_LOOP_3_quantized_value_slc_63_32_cse_slc , (APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm[55:39])})
      + 26'b00000000000000000000000001;
  assign QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_nl = nl_QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_nl[25:0];
  assign QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1 = readslicef_26_1_25(QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_nl);
  assign attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0_mx0w6 = MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0, or_dcpl_1145);
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48_mx0w2 = MUX_v_24_16_2(attention_2_1_16_16_4_4_k_proj_re_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_1_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_3_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_4_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_5_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_6_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_7_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_8_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_9_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_10_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_11_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_12_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_13_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_14_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_15_sva_1_39_16, {reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2});
  assign attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16_mx0w5 = MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1,
      attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16, or_dcpl_1145);
  assign attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16, or_dcpl_1085);
  assign attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16, or_dcpl_1083);
  assign attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16, or_dcpl_1071);
  assign attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16, or_dcpl_1073);
  assign attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16, or_dcpl_1091);
  assign attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16, or_dcpl_1090);
  assign attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16, or_dcpl_1089);
  assign attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16, or_dcpl_1088);
  assign attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16, or_dcpl_1087);
  assign attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16, or_dcpl_1086);
  assign attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1,
      attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16, or_dcpl_1067);
  assign attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16, or_dcpl_1152);
  assign attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16, or_dcpl_1155);
  assign attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16, or_dcpl_1156);
  assign attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16, or_dcpl_1158);
  assign attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16, or_dcpl_1159);
  assign attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16, or_dcpl_1160);
  assign attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16, or_dcpl_1161);
  assign attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16, or_dcpl_1162);
  assign attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16, or_dcpl_1164);
  assign attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16, or_dcpl_1165);
  assign attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16, or_dcpl_1166);
  assign attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16, or_dcpl_1167);
  assign attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16, or_dcpl_1168);
  assign attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16, or_dcpl_1169);
  assign attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1,
      attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16, or_dcpl_1170);
  assign attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16, or_dcpl_1133);
  assign attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16, or_dcpl_1108);
  assign attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16, or_dcpl_1132);
  assign attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16, or_dcpl_1114);
  assign attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16, or_dcpl_1131);
  assign attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16, or_dcpl_1116);
  assign attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16, or_dcpl_1130);
  assign attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16, or_dcpl_1118);
  assign attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16, or_dcpl_1128);
  assign attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16, or_dcpl_1120);
  assign attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16, or_dcpl_1127);
  assign attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16, or_dcpl_1121);
  assign attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16, or_dcpl_1126);
  assign attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16, or_dcpl_1122);
  assign attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16, or_dcpl_1125);
  assign attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1,
      attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16, or_dcpl_1123);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_7 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7, attention_2_1_16_16_4_4_quantized_hidden_states_0_6_sva_7,
      attention_2_1_16_16_4_4_quantized_hidden_states_0_7_sva_7, attention_2_1_16_16_4_4_quantized_hidden_states_0_8_sva_7,
      attention_2_1_16_16_4_4_quantized_hidden_states_0_9_sva_7, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_7, {reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_6 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_1,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_6, {reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_5 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_2,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_5, {reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_4 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_3,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_4, {reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_3 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_4,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_3, {reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_2 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_5,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_2, {reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_1 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_6,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_1, {reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_0 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_7,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_0, {reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_7 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7, attention_2_1_16_16_4_4_quantized_hidden_states_0_6_sva_7,
      attention_2_1_16_16_4_4_quantized_hidden_states_0_7_sva_7, attention_2_1_16_16_4_4_quantized_hidden_states_0_8_sva_7,
      attention_2_1_16_16_4_4_quantized_hidden_states_0_9_sva_7, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_7, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_6 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_1,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_6, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_5 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_2,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_5, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_4 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_3,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_4, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_3 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_4,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_3, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_2 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_5,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_2, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_1 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_6,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_1, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_0 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_7,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_0, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_7 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7, attention_2_1_16_16_4_4_quantized_hidden_states_0_6_sva_7,
      attention_2_1_16_16_4_4_quantized_hidden_states_0_7_sva_7, attention_2_1_16_16_4_4_quantized_hidden_states_0_8_sva_7,
      attention_2_1_16_16_4_4_quantized_hidden_states_0_9_sva_7, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_7, {reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_6 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_1,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_6, {reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_5 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_2,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_5, {reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_4 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_3,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_4, {reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_3 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_4,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_3, {reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_2 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_5,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_2, {reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_1 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_6,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_1, {reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_0 = MUX_s_1_16_2(reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_7,
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse, reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse,
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse, attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0, attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0, attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0,
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_0, {reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign nl_LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_2 = conv_u2s_2_3({LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1
      , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0}) + 3'b001;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_2 = nl_LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_2[2:0];
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm = (LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_0
      & (~ LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_1))
      | LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1;
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux_32_nl = MUX_v_24_16_2(attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16, attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16, attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16, attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16, attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16, attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16, attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16, attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16, {reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_7,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_7), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_nl = LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_1_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_6,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_6), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_3_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_1_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_2_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_5,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_5), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_4_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_2_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_3_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_4,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_4), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_5_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_3_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_4_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_3,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_3), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_6_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_4_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_5_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_2,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_2), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_7_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_5_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_6_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_1,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_1), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_8_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_6_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_7_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_0,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_2_new_val_sva_3_0), LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_9_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_2_mux_7_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_2_or_itm;
  assign nl_operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1 = operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux_32_nl
      + conv_s2s_8_24({LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_nl
      , LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_3_nl ,
      LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_4_nl , LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_5_nl
      , LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_6_nl ,
      LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_7_nl , LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_8_nl
      , LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_9_nl});
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1 = nl_operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_acc_psp_sva_1[23:0];
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_LINEAR_FORWARD_NO_MUL_LOOP_4_2_and_1_cse_1
      = LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_1
      & (~ LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_0);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_1
      = MUX_s_1_4_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7,
      {reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_2_weight_val_conc_1_1_1_0_svs_1_0
      = MUX_s_1_4_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6,
      {reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_17_nl = MUX_v_24_16_2(attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16, attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16, attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16, attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16, attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16, attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16, attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16, attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16, {reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_7,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_7), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_nl = LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_1_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_6,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_6), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_5_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_1_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_2_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_5,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_5), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_6_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_2_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_3_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_4,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_4), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_7_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_3_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_4_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_3,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_3), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_8_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_4_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_5_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_2,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_2), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_9_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_5_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_6_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_1,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_10_nl
      = LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_6_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_7_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_0,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_1_new_val_sva_3_0), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_11_nl
      = LINEAR_FORWARD_NO_MUL_LOOP_4_1_mux_7_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign nl_operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1 = operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_17_nl
      + conv_s2s_8_24({LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_nl
      , LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_5_nl ,
      LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_6_nl , LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_7_nl
      , LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_8_nl ,
      LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_9_nl , LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_10_nl
      , LINEAR_FORWARD_NO_MUL_LOOP_4_1_LINEAR_FORWARD_NO_MUL_LOOP_4_1_and_11_nl});
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1 = nl_operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_acc_psp_sva_1[23:0];
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1
      = (LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_conc_1_1_1_0_svs_1==2'b10);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_conc_1_1_1_0_svs_1
      = MUX_v_2_4_2((reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3[1:0]),
      (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3[3:2]),
      (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3[5:4]),
      (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3[7:6]),
      {reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm = (LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_0
      & (~ LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_1))
      | LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1;
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_17_nl = MUX_v_24_16_2(attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16, attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16, attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16, attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16, attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16, attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16, attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16, attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16, {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
      , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_mux_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_7,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_7), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_nl = LINEAR_FORWARD_NO_MUL_LOOP_4_mux_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_mux_1_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_6,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_6), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_3_nl = LINEAR_FORWARD_NO_MUL_LOOP_4_mux_1_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_mux_2_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_5,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_5), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_4_nl = LINEAR_FORWARD_NO_MUL_LOOP_4_mux_2_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_mux_3_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_4,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_4), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_5_nl = LINEAR_FORWARD_NO_MUL_LOOP_4_mux_3_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_mux_4_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_3,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_3), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_6_nl = LINEAR_FORWARD_NO_MUL_LOOP_4_mux_4_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_mux_5_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_2,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_2), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_7_nl = LINEAR_FORWARD_NO_MUL_LOOP_4_mux_5_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_mux_6_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_1,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_1), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_8_nl = LINEAR_FORWARD_NO_MUL_LOOP_4_mux_6_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_mux_7_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_0,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_new_val_sva_3_0), LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_9_nl = LINEAR_FORWARD_NO_MUL_LOOP_4_mux_7_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_or_itm;
  assign nl_operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1 = operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_17_nl
      + conv_s2s_8_24({LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_nl
      , LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_3_nl , LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_4_nl
      , LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_5_nl , LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_6_nl
      , LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_7_nl , LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_8_nl
      , LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_9_nl});
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1 = nl_operator_40_24_true_AC_TRN_AC_WRAP_8_true_acc_psp_sva_1[23:0];
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_LINEAR_FORWARD_NO_MUL_LOOP_4_and_1_cse_1 =
      LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_1
      & (~ LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_0);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_1
      = MUX_s_1_4_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7,
      {LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1 , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_weight_val_conc_1_1_1_0_svs_1_0
      = MUX_s_1_4_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4, reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6,
      {LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1 , LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0});
  assign RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1
      = MUX_v_24_16_2(attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16,
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_39_16, apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_3_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_re_0_7_sva_2_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_3_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16,
      attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_3_39_16,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1});
  assign GEMM_3D_FLOAT_LOOP_3_and_tmp_4_sva_mx0w2 = GEMM_3D_FLOAT_LOOP_3_and_stg_1_3_sva_1
      & (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2:1]==2'b01);
  assign GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_0_sva_mx0w3 = nor_1229_cse & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign GEMM_3D_FLOAT_LOOP_3_and_tmp_5_sva_mx0w2 = GEMM_3D_FLOAT_LOOP_3_and_stg_1_2_sva_1
      & (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2:1]==2'b01);
  assign GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_1_sva_mx0w3 = GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_1_sva_1
      & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign GEMM_3D_FLOAT_LOOP_3_and_tmp_6_sva_mx0w1 = GEMM_3D_FLOAT_LOOP_3_and_stg_1_1_sva_1
      & (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2:1]==2'b01);
  assign GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva_mx0w3 = GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_2_sva_1
      & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign GEMM_3D_FLOAT_LOOP_3_and_tmp_7_sva_mx0w1 = GEMM_3D_FLOAT_LOOP_3_and_stg_1_0_sva_1
      & (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2:1]==2'b01);
  assign GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva_mx0w3 = GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_3_sva_1
      & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1
      = MUX_v_24_8_2(attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_39_16, attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8
      = MUX_v_8_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[15:8]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_8,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_15_8, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[15:8]),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[15:8]), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[15:8]),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[15:8]), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[15:8]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[7]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_7,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_7, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[7]),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[7]), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[7]),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[7]), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[7]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[6]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_6,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_6, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[6]),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[6]), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[6]),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[6]), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[6]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[5]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_5,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_5, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[5]),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[5]), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[5]),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[5]), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[5]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[4]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_4,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_4, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[4]),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[4]), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[4]),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[4]), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[4]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[3]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_3,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_3, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[3]),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[3]), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[3]),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[3]), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[3]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[2]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_2,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_2, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[2]),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[2]), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[2]),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[2]), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[2]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[1]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_1,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_1, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[1]),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[1]), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[1]),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[1]), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[1]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[0]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_0,
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_0, (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[0]),
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[0]), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[0]),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[0]), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[0]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1
      = MUX_v_24_8_2(attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_39_16, attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_39_16,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm
      = MUX_v_8_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[15:8]), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[15:8]),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[7]), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[7]),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_7, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_7, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_7, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_7,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[6]), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[6]),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_6, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_6, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_6, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_6,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[5]), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[5]),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_5, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_5, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_5, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_5,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[4]), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[4]),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_4, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_4, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_4, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_4,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[3]), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[3]),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_3, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_3, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_3, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_3,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[2]), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[2]),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_2, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_2, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_2, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_2,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[1]), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[1]),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_1, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_1, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_1, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_1,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[0]), (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[0]),
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_0, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_0, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_0, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_0,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_1_nl
      = MUX_v_24_8_2(attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_7_nl
      = MUX_v_8_8_2(attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_8, reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_ftd,
      ({attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_13 , (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[12:8])}),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_8, (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0[15:8]),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0[15:8]), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0[15:8]),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0[15:8]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_25_nl
      = MUX_v_8_8_2(({reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd ,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_1 , reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_2
      , reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_3 , reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_4
      , reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_5 , reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_6
      , reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_7}), ({reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd
      , reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_1 , reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_2
      , reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_3 , reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_4
      , reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_5 , reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_6
      , reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_7}), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[7:0]),
      ({attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_7 , attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_6
      , attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_5 , attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_4
      , attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_3 , attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_2
      , attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_1 , attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_0}),
      (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0[7:0]), (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0[7:0]),
      (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0[7:0]), (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0[7:0]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign nl_APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1 = ({(~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_1_nl)
      , (~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_7_nl)
      , (~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_25_nl)})
      + 40'b0000000000000000000000000000000000000001;
  assign APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1 = nl_APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1[39:0];
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_nl
      = MUX_v_24_8_2(attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_39_16,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_6_nl
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[15]), attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_15,
      (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8[7]), (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8[7]),
      (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8[7]), (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8[7]),
      (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8[7]), (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8[7]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_26_nl
      = MUX_v_3_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[14:12]), attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_14_12,
      (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8[6:4]), (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8[6:4]),
      (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8[6:4]), (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8[6:4]),
      (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8[6:4]), (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8[6:4]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_27_nl
      = MUX_v_3_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[11:9]), attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_11_9,
      (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8[3:1]), (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8[3:1]),
      (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8[3:1]), (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8[3:1]),
      (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8[3:1]), (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8[3:1]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_28_nl
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[8]), attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_8,
      (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8[0]), (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8[0]),
      (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8[0]), (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8[0]),
      (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8[0]), (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8[0]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_16_nl
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[7]), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[7]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_7, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_7, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_7, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_7,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_17_nl
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[6]), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[6]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_6, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_6, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_6, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_6,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_18_nl
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[5]), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[5]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_5, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_5, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_5, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_5,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_19_nl
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[4]), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[4]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_4, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_4, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_4, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_4,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_20_nl
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[3]), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[3]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_3, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_3, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_3, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_3,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_21_nl
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[2]), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[2]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_2, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_2, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_2, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_2,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_22_nl
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[1]), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[1]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_1, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_1, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_1, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_1,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_23_nl
      = MUX_s_1_8_2((attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[0]), (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[0]),
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_0, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_0, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_0, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_0,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign nl_APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1 = ({(~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_nl)
      , (~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_6_nl)
      , (~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_26_nl)
      , (~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_27_nl)
      , (~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_28_nl)
      , (~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_16_nl)
      , (~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_17_nl)
      , (~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_18_nl)
      , (~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_19_nl)
      , (~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_20_nl)
      , (~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_21_nl)
      , (~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_22_nl)
      , (~ APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_23_nl)})
      + 40'b0000000000000000000000000000000000000001;
  assign APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1 = nl_APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1[39:0];
  assign RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_39_16_1
      = MUX_v_24_16_2(attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_39_16, attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_39_16,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1});
  assign RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1
      = MUX_v_16_16_2(attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_15_0, ({attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_15_8
      , attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_7 , attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_6
      , attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_5 , attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_4
      , attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_3 , attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_2
      , attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_1 , attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_0}),
      attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_15_0, attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_15_0,
      attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_15_0, attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_15_0,
      attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_15_0, attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_15_0,
      attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_15_0, attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_15_0,
      ({attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_15_13 , attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0}),
      ({attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_15_8 , attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_7
      , attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_6 , attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_5
      , attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_4 , attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_3
      , attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_2 , attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_1
      , attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_0}), attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_15_0,
      attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_15_0, attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_15_0,
      attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_15_0, {reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1});
  assign attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx1 = MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_3,
      CM_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_ctmp_sva_1, CM_LOOP_3_acc_tmp[2]);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx2 = MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z[39:0]),
      attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_4, or_dcpl_1178);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx1 = MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z[39:0]),
      attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_5, or_dcpl_1180);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx1 = MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z[39:0]),
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_5, or_dcpl_1181);
  assign nand_378_nl = ~(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 & (CM_LOOP_3_acc_tmp[0]));
  assign attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx1 = MUX_v_40_2_2(CM_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_ctmp_sva_1,
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_3, nand_378_nl);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx2 = MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z[39:0]),
      attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_4, or_dcpl_1183);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx1 = MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z[39:0]),
      attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_4, or_dcpl_1184);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx1 = MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z[39:0]),
      attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_4, or_dcpl_1186);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx1 = MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z[39:0]),
      attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_4, or_dcpl_1187);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx1 = MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_3,
      CM_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_ctmp_sva_1, CM_LOOP_3_acc_tmp[1]);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx2 = MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z[39:0]),
      attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_4, or_dcpl_1188);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx1 = MUX_v_40_2_2((SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z[39:0]),
      attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_4, or_dcpl_1189);
  assign nl_APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_nl = APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm
      + APPLY_ROTARY_POS_EMB_LOOP_6_mul_3_itm;
  assign APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_nl = nl_APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_nl[55:0];
  assign APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1 = readslicef_56_40_16(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_nl);
  assign nl_APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_nl = APPLY_ROTARY_POS_EMB_LOOP_6_mul_itm
      + APPLY_ROTARY_POS_EMB_LOOP_6_mul_1_itm;
  assign APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_nl = nl_APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_nl[55:0];
  assign APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1 = readslicef_56_40_16(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_nl);
  assign nl_CACHE_UPDATE_LOOP_3_acc_sdt_1 = conv_u2u_2_3({reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1}) + conv_u2u_2_3(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2);
  assign CACHE_UPDATE_LOOP_3_acc_sdt_1 = nl_CACHE_UPDATE_LOOP_3_acc_sdt_1[2:0];
  assign nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_15_sdt_1 = conv_u2u_2_3(TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3[2:1])
      + conv_u2u_2_3({reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_15_sdt_1 = nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_15_sdt_1[2:0];
  assign nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_sdt_1 = conv_u2u_2_3({reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1}) + conv_u2u_2_3({reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_sdt_1 = nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_sdt_1[2:0];
  assign GEMM_3D_FLOAT_LOOP_3_and_tmp_sva_mx0w0 = GEMM_3D_FLOAT_LOOP_3_and_stg_2_3_sva_1
      & (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2]);
  assign GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva_mx0w0 = GEMM_3D_FLOAT_LOOP_3_and_stg_2_0_sva_1
      & (~ (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2]));
  assign GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva_mx0w0 = GEMM_3D_FLOAT_LOOP_3_and_stg_2_2_sva_1
      & (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2]);
  assign GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva_mx0w0 = GEMM_3D_FLOAT_LOOP_3_and_stg_2_1_sva_1
      & (~ (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2]));
  assign GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva_mx0w0 = GEMM_3D_FLOAT_LOOP_3_and_stg_2_1_sva_1
      & (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2]);
  assign GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva_mx0w0 = GEMM_3D_FLOAT_LOOP_3_and_stg_2_2_sva_1
      & (~ (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2]));
  assign GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva_mx0w0 = GEMM_3D_FLOAT_LOOP_3_and_stg_2_0_sva_1
      & (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2]);
  assign GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva_mx0w0 = GEMM_3D_FLOAT_LOOP_3_and_stg_2_3_sva_1
      & (~ (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2]));
  assign GEMM_3D_FLOAT_LOOP_3_and_stg_2_0_sva_1 = GEMM_3D_FLOAT_LOOP_3_and_stg_1_0_sva_1
      & (~ (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[1]));
  assign GEMM_3D_FLOAT_LOOP_3_and_stg_2_1_sva_1 = GEMM_3D_FLOAT_LOOP_3_and_stg_1_1_sva_1
      & (~ (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[1]));
  assign GEMM_3D_FLOAT_LOOP_3_and_stg_2_2_sva_1 = GEMM_3D_FLOAT_LOOP_3_and_stg_1_2_sva_1
      & (~ (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[1]));
  assign GEMM_3D_FLOAT_LOOP_3_and_stg_2_3_sva_1 = GEMM_3D_FLOAT_LOOP_3_and_stg_1_3_sva_1
      & (~ (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[1]));
  assign GEMM_3D_FLOAT_LOOP_3_and_stg_1_0_sva_1 = ~((z_out_11[0]) | (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[0]));
  assign GEMM_3D_FLOAT_LOOP_3_and_stg_1_1_sva_1 = (z_out_11[0]) & (~ (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[0]));
  assign GEMM_3D_FLOAT_LOOP_3_and_stg_1_2_sva_1 = (~ (z_out_11[0])) & (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[0]);
  assign GEMM_3D_FLOAT_LOOP_3_and_stg_1_3_sva_1 = (z_out_11[0]) & (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[0]);
  assign nl_GEMM_3D_FLOAT_LOOP_4_acc_sdt_1 = conv_u2u_2_3(GEMM_3D_FLOAT_LOOP_4_acc_13_sdt_1[2:1])
      + conv_u2u_2_3({reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign GEMM_3D_FLOAT_LOOP_4_acc_sdt_1 = nl_GEMM_3D_FLOAT_LOOP_4_acc_sdt_1[2:0];
  assign nl_GEMM_3D_FLOAT_LOOP_4_acc_13_sdt_1 = conv_u2u_2_3(z_out_11[2:1]) + conv_u2u_2_3({reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign GEMM_3D_FLOAT_LOOP_4_acc_13_sdt_1 = nl_GEMM_3D_FLOAT_LOOP_4_acc_13_sdt_1[2:0];
  assign or_3014_nl = or_dcpl_1196 | or_dcpl_1195;
  assign attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6_mx1 = MUX_v_40_2_2(({{1{SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1[38]}},
      SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1}), attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6,
      or_3014_nl);
  assign or_3017_nl = or_dcpl_1199 | or_dcpl_1198;
  assign attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6_mx1 = MUX_v_40_2_2(({{1{SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1[38]}},
      SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1}), attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6,
      or_3017_nl);
  assign or_3019_nl = or_dcpl_1196 | or_dcpl_1201;
  assign attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6_mx1 = MUX_v_40_2_2(({{1{SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1[38]}},
      SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1}), attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6,
      or_3019_nl);
  assign or_3021_nl = or_dcpl_1199 | or_dcpl_1203;
  assign attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6_mx1 = MUX_v_40_2_2(({{1{SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1[38]}},
      SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1}), attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6,
      or_3021_nl);
  assign or_3022_nl = or_dcpl_1196 | or_dcpl_1203;
  assign attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6_mx1 = MUX_v_40_2_2(({{1{SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1[38]}},
      SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1}), attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6,
      or_3022_nl);
  assign or_3023_nl = or_dcpl_1199 | or_dcpl_1201;
  assign attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6_mx1 = MUX_v_40_2_2(({{1{SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1[38]}},
      SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1}), attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6,
      or_3023_nl);
  assign or_3024_nl = or_dcpl_1196 | or_dcpl_1198;
  assign attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6_mx1 = MUX_v_40_2_2(({{1{SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1[38]}},
      SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1}), attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6,
      or_3024_nl);
  assign or_3025_nl = or_dcpl_1199 | or_dcpl_1195;
  assign attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6_mx1 = MUX_v_40_2_2(({{1{SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1[38]}},
      SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1}), attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6,
      or_3025_nl);
  assign or_3027_nl = or_dcpl_1209 | or_dcpl_1195;
  assign attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6_mx1 = MUX_v_40_2_2(({{1{SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1[38]}},
      SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1}), attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6,
      or_3027_nl);
  assign or_3028_nl = or_dcpl_1209 | or_dcpl_1198;
  assign attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6_mx1 = MUX_v_40_2_2(({{1{SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1[38]}},
      SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1}), attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6,
      or_3028_nl);
  assign or_3029_nl = or_dcpl_1209 | or_dcpl_1201;
  assign attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6_mx1 = MUX_v_40_2_2(({{1{SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1[38]}},
      SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1}), attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6,
      or_3029_nl);
  assign or_3030_nl = or_dcpl_1209 | or_dcpl_1203;
  assign attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6_mx1 = MUX_v_40_2_2(({{1{SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1[38]}},
      SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1}), attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6,
      or_3030_nl);
  assign SF_LOOP_3_and_nl = (SF_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_psp_sva_1[39])
      & (SF_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_psp_sva_1[0]);
  assign nl_SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1 = (SF_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_psp_sva_1[39:1])
      + conv_u2s_1_39(SF_LOOP_3_and_nl);
  assign SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1 = nl_SF_LOOP_3_SF_LOOP_3_SF_LOOP_3_acc_psp_sva_1[38:0];
  assign SF_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_psp_sva_1 = MUX_v_40_12_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6,
      attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6, attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6,
      attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6, attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6,
      attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6, attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6,
      attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6, attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6,
      attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6, attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6,
      attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign CM_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_ctmp_sva_1 =
      MUX_v_40_4_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_3, attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_3,
      attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_3, attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_3,
      {reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign nl_CM_LOOP_3_acc_tmp = conv_u2u_1_3(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd)
      + conv_u2u_2_3({reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign CM_LOOP_3_acc_tmp = nl_CM_LOOP_3_acc_tmp[2:0];
  assign attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8_mx1 = MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8, or_dcpl_1178);
  assign attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9_mx1 = MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9, or_dcpl_1063);
  assign attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8_mx1 = MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8, or_dcpl_1187);
  assign attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8_mx1 = MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8, or_dcpl_1183);
  assign attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9_mx1 = MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9, or_dcpl_1181);
  assign attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8_mx1 = MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8, or_dcpl_1188);
  assign attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8_mx1 = MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8, or_dcpl_1081);
  assign attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9_mx1 = MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9, or_dcpl_1076);
  assign attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8_mx1 = MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8, or_dcpl_1186);
  assign attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8_mx1 = MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8, or_dcpl_1184);
  assign attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9_mx1 = MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9, or_dcpl_1180);
  assign attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8_mx1 = MUX_v_40_2_2(SOFTMAX_LOOP_4_acc_3_cse_sva_1,
      attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8, or_dcpl_1189);
  assign SOFTMAX_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_cse_sva_1
      = MUX_v_40_15_2(attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1, attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_3,
      attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_3, attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1, attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_3,
      attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_3, attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1, attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_3,
      attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_3, attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1, attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_3,
      attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_3, {reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign nl_operator_40_24_true_AC_TRN_AC_WRAP_acc_nl = ({operator_80_48_true_AC_TRN_AC_WRAP_operator_80_48_true_AC_TRN_AC_WRAP_slc_SOFTMAX_LOOP_4_sqr_56_1_itm_slc
      , (APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm[55:33])}) + 24'b000000000000000000000001;
  assign operator_40_24_true_AC_TRN_AC_WRAP_acc_nl = nl_operator_40_24_true_AC_TRN_AC_WRAP_acc_nl[23:0];
  assign nl_SOFTMAX_LOOP_4_acc_3_cse_sva_1 = ({operator_40_24_true_AC_TRN_AC_WRAP_acc_nl
      , (APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm[32:17])}) + GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm;
  assign SOFTMAX_LOOP_4_acc_3_cse_sva_1 = nl_SOFTMAX_LOOP_4_acc_3_cse_sva_1[39:0];
  assign GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva_mx0w0 = GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_3_sva_1
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva_mx0w0 = GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_2_sva_1
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva_mx0w0 = GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_1_sva_1
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva_mx0w0 = nor_1229_cse & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_1_sva_1 = reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd);
  assign GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_2_sva_1 = (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1)
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd;
  assign GEMM_3D_FLOAT_LOOP_3_1_and_stg_1_3_sva_1 = reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd;
  assign nl_GEMM_3D_FLOAT_LOOP_4_1_acc_12_sdt_1 = conv_u2u_2_3({reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1}) + conv_u2u_2_3(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2);
  assign GEMM_3D_FLOAT_LOOP_4_1_acc_12_sdt_1 = nl_GEMM_3D_FLOAT_LOOP_4_1_acc_12_sdt_1[2:0];
  assign nl_attention_abs_5_qr_sva_1 = conv_u2s_39_40(~ (attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_2_mx0[38:0]))
      + 40'b0000000000000000000000000000000000000001;
  assign attention_abs_5_qr_sva_1 = nl_attention_abs_5_qr_sva_1[39:0];
  assign attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_2_mx0 = MUX_v_40_2_2(RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1, or_dcpl_1108);
  assign nl_attention_abs_6_mux_2 = conv_u2s_39_40(~ (RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva[38:0]))
      + 40'b0000000000000000000000000000000000000001;
  assign attention_abs_6_mux_2 = nl_attention_abs_6_mux_2[39:0];
  assign QUANTIZE_ACTIVATION_LOOP_2_1_attention_abs_6_nand_nl = ~((attention_abs_6_mux_2[39])
      & (RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva[39]));
  assign attention_abs_6_mux_3_nl = MUX_v_39_2_2((RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva[38:0]),
      (attention_abs_6_mux_2[38:0]), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva[39]);
  assign nl_QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_nl = conv_s2u_40_41({reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      , QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_38_0}) + conv_s2u_40_41({QUANTIZE_ACTIVATION_LOOP_2_1_attention_abs_6_nand_nl
      , (~ attention_abs_6_mux_3_nl)}) + 41'b00000000000000000000000000000000000000001;
  assign QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_nl = nl_QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_nl[40:0];
  assign QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_itm_40_1 = readslicef_41_1_40(QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_nl);
  assign RMS_NORM_LOOP_2_2_and_29_ssc_1 = (~ QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_itm_40_1)
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign RMS_NORM_LOOP_2_2_and_34_ssc_1 = (RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva[39])
      & RMS_NORM_LOOP_2_2_and_30_m1c_1;
  assign RMS_NORM_LOOP_2_2_and_30_m1c_1 = QUANTIZE_ACTIVATION_LOOP_2_1_acc_4_itm_40_1
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_nor_1_ssc_1 = ~((attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1[39])
      | reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign RMS_NORM_LOOP_2_2_and_33_ssc_1 = (~ (RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva[39]))
      & RMS_NORM_LOOP_2_2_and_30_m1c;
  assign nl_QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_nl = ({1'b1
      , reg_QUANTIZE_ACTIVATION_LOOP_3_quantized_value_slc_63_32_cse_slc , (APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm[55:39])})
      + 26'b00000000000000000000000001;
  assign QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_nl = nl_QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_nl[25:0];
  assign QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1 = readslicef_26_1_25(QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_nl);
  assign QUANTIZE_ACTIVATION_LOOP_3_1_nand_seb_1 = ~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2==2'b11) & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd);
  assign output_0_15_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_15_lpi_4_39_16, or_dcpl_1152);
  assign output_0_0_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_0_lpi_4_39_16, or_dcpl_1155);
  assign output_0_14_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_14_lpi_4_39_16, or_dcpl_1156);
  assign output_0_1_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_1_lpi_4_39_16, or_dcpl_1158);
  assign output_0_13_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_13_lpi_4_39_16, or_dcpl_1159);
  assign output_0_2_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_2_lpi_4_39_16, or_dcpl_1160);
  assign output_0_12_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_12_lpi_4_39_16, or_dcpl_1161);
  assign output_0_3_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_3_lpi_4_39_16, or_dcpl_1162);
  assign output_0_11_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_11_lpi_4_39_16, or_dcpl_1164);
  assign output_0_4_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_4_lpi_4_39_16, or_dcpl_1165);
  assign output_0_10_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_10_lpi_4_39_16, or_dcpl_1166);
  assign output_0_5_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_5_lpi_4_39_16, or_dcpl_1167);
  assign output_0_9_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_9_lpi_4_39_16, or_dcpl_1168);
  assign output_0_6_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_6_lpi_4_39_16, or_dcpl_1169);
  assign output_0_8_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_8_lpi_4_39_16, or_dcpl_1170);
  assign output_0_7_lpi_4_39_16_mx1 = MUX_v_24_2_2(operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1,
      output_0_7_lpi_4_39_16, or_dcpl_1141);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_7_1 = MUX_s_1_16_2(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva,
      attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_7, attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_7,
      attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_7, attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_7,
      attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_7, attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_7,
      attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_7, attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_7,
      attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_7, attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_7,
      attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_7, attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_7,
      attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_7, attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_7,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_7, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_0_1 = MUX_s_1_16_2(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_6_1 = MUX_s_1_16_2(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_1_1 = MUX_s_1_16_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_5_1 = MUX_s_1_16_2(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_2_1 = MUX_s_1_16_2(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_4_1 = MUX_s_1_16_2(LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_3_1 = MUX_s_1_16_2(reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse,
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse, reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse,
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_mux_32_nl = MUX_v_24_16_2(output_0_0_lpi_4_39_16,
      output_0_1_lpi_4_39_16, output_0_2_lpi_4_39_16, output_0_3_lpi_4_39_16, output_0_4_lpi_4_39_16,
      output_0_5_lpi_4_39_16, output_0_6_lpi_4_39_16, output_0_7_lpi_4_39_16, output_0_8_lpi_4_39_16,
      output_0_9_lpi_4_39_16, output_0_10_lpi_4_39_16, output_0_11_lpi_4_39_16, output_0_12_lpi_4_39_16,
      output_0_13_lpi_4_39_16, output_0_14_lpi_4_39_16, output_0_15_lpi_4_39_16,
      {reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2});
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_7_1,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_7_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_nl = LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_nl
      & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_1_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_6_1,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_6_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_3_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_1_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_2_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_5_1,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_5_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_4_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_2_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_3_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_4_1,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_4_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_5_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_3_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_4_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_3_1,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_3_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_6_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_4_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_5_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_2_1,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_2_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_7_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_5_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_6_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_1_1,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_1_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_8_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_6_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_7_nl = MUX_s_1_2_2(LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_0_1,
      (~ LINEAR_FORWARD_NO_MUL_LOOP_4_3_new_val_sva_1_0_1), LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_9_nl =
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_mux_7_nl & LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0;
  assign nl_operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1 = operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_mux_32_nl
      + conv_s2s_8_24({LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_nl
      , LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_3_nl ,
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_4_nl , LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_5_nl
      , LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_6_nl ,
      LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_7_nl , LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_8_nl
      , LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_9_nl});
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1 = nl_operator_40_24_true_AC_TRN_AC_WRAP_8_true_3_acc_psp_sva_1[23:0];
  assign nl_CACHE_UPDATE_LOOP_2_1_acc_2_nl = ({1'b1 , (z_out_4[1:0])}) + 3'b001;
  assign CACHE_UPDATE_LOOP_2_1_acc_2_nl = nl_CACHE_UPDATE_LOOP_2_1_acc_2_nl[2:0];
  assign CACHE_UPDATE_LOOP_2_1_acc_2_itm_2_1 = readslicef_3_1_2(CACHE_UPDATE_LOOP_2_1_acc_2_nl);
  assign nl_attention_max_attn_fixed_t_1_acc_1_nl = conv_s2u_40_41({(~ reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1)
      , (~ reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1)}) + 41'b00000000000000000000000000000000000000001;
  assign attention_max_attn_fixed_t_1_acc_1_nl = nl_attention_max_attn_fixed_t_1_acc_1_nl[40:0];
  assign attention_max_attn_fixed_t_1_acc_1_itm_40_1 = readslicef_41_1_40(attention_max_attn_fixed_t_1_acc_1_nl);
  assign LINEAR_FORWARD_NO_MUL_LOOP_4_1_exs_2_0 = ((LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_slc_LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_LINEAR_FORWARD_NO_MUL_LOOP_4_3_weight_val_conc_1_1_1_0_svs_1==2'b01))
      | LINEAR_FORWARD_NO_MUL_LOOP_4_3_LINEAR_FORWARD_NO_MUL_LOOP_4_3_and_1_cse_1;
  assign nl_CACHE_UPDATE_LOOP_2_acc_2_nl = ({1'b1 , (z_out_3[1:0])}) + 3'b001;
  assign CACHE_UPDATE_LOOP_2_acc_2_nl = nl_CACHE_UPDATE_LOOP_2_acc_2_nl[2:0];
  assign CACHE_UPDATE_LOOP_2_acc_2_itm_2_1 = readslicef_3_1_2(CACHE_UPDATE_LOOP_2_acc_2_nl);
  assign nl_SOFTMAX_LOOP_3_acc_3_nl = conv_s2u_40_41({QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39
      , QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0}) - conv_s2u_40_41(SOFTMAX_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_cse_sva_1);
  assign SOFTMAX_LOOP_3_acc_3_nl = nl_SOFTMAX_LOOP_3_acc_3_nl[40:0];
  assign SOFTMAX_LOOP_3_acc_3_itm_40_1 = readslicef_41_1_40(SOFTMAX_LOOP_3_acc_3_nl);
  assign CACHE_UPDATE_LOOP_1_and_tmp = (z_out_3[2]) & (z_out_5[2]);
  assign RESHAPE_2D_TO_3D_LOOP_2_2_and_cse = (z_out_5[2]) & (z_out_4[2]);
  assign for_for_and_tmp = (LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1[4]) & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4;
  assign or_dcpl_4 = reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd | (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign and_dcpl = ~((fsm_output[3]) | (fsm_output[6]));
  assign and_dcpl_1 = ~((fsm_output[8]) | (fsm_output[5]));
  assign or_tmp_11 = (fsm_output[2]) | (~ (fsm_output[4]));
  assign nor_646_cse = ~((fsm_output[5:4]!=2'b00));
  assign or_tmp_48 = (~ (fsm_output[4])) | (fsm_output[8]);
  assign or_dcpl_45 = ~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]) & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  assign or_dcpl_47 = ~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]==2'b11));
  assign or_dcpl_54 = ~(reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign or_dcpl_60 = (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0])) | reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1;
  assign or_133_cse = (fsm_output[4]) | (fsm_output[8]);
  assign or_dcpl_68 = (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]) | (~ reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  assign or_dcpl_79 = (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]) | reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1;
  assign or_dcpl_96 = (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd) | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign or_241_cse = (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b00);
  assign or_tmp_104 = (fsm_output[1]) | (fsm_output[8]);
  assign or_255_cse = (fsm_output[4]) | (fsm_output[2]);
  assign or_262_cse = (~ (fsm_output[1])) | (fsm_output[8]);
  assign mux_tmp_87 = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), fsm_output[2]);
  assign mux_tmp_91 = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), fsm_output[5]);
  assign nor_tmp_28 = (fsm_output[6]) & (fsm_output[8]);
  assign mux_tmp_121 = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), fsm_output[6]);
  assign and_dcpl_26 = ~((fsm_output[8:7]!=2'b00));
  assign or_349_cse = (fsm_output[1]) | (fsm_output[0]) | (fsm_output[2]) | (fsm_output[5])
      | (fsm_output[4]);
  assign nand_129_cse = ~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd);
  assign or_361_cse = (fsm_output[8:7]!=2'b01);
  assign or_362_cse = (fsm_output[8:7]!=2'b00);
  assign mux_304_cse = MUX_s_1_2_2(or_361_cse, or_362_cse, fsm_output[6]);
  assign and_dcpl_45 = (fsm_output[7:6]==2'b10);
  assign nor_tmp_99 = (fsm_output[4]) & (fsm_output[8]);
  assign and_dcpl_57 = (fsm_output[7:6]==2'b01);
  assign and_dcpl_61 = ~((fsm_output[8]) | (fsm_output[4]));
  assign or_619_cse = (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd) |
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1]);
  assign and_dcpl_65 = (fsm_output[1]) & (fsm_output[3]);
  assign or_dcpl_332 = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b00);
  assign or_dcpl_337 = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b10);
  assign or_dcpl_342 = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b01);
  assign or_dcpl_351 = ~((reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2==2'b11));
  assign or_dcpl_377 = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd;
  assign or_750_cse = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0])
      | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  assign or_753_cse = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0])
      | (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  assign or_tmp_330 = ~((fsm_output[1]) & (fsm_output[0]) & (fsm_output[2]) & (~
      (fsm_output[4])));
  assign or_790_cse = (~ (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0]))
      | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  assign nand_143_cse = ~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd &
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1]));
  assign or_806_cse = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd | (~ (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1]));
  assign or_822_cse = (fsm_output[8:7]!=2'b10);
  assign nor_tmp_117 = or_1984_cse & (fsm_output[8]);
  assign mux_tmp_363 = MUX_s_1_2_2((fsm_output[7]), (fsm_output[8]), fsm_output[6]);
  assign not_tmp_253 = ~((fsm_output[6:4]==3'b111));
  assign or_dcpl_508 = (~ reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd) | reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1;
  assign or_dcpl_512 = ~(reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd & reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1);
  assign or_dcpl_584 = reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign or_tmp_464 = (~ (fsm_output[6])) | (fsm_output[8]);
  assign nor_717_cse = ~((fsm_output[2:1]!=2'b00));
  assign mux_528_cse = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), fsm_output[4]);
  assign or_dcpl_672 = (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b10);
  assign or_tmp_507 = (fsm_output[8:6]!=3'b011);
  assign or_1197_cse = (fsm_output[8:6]!=3'b100);
  assign mux_tmp_604 = MUX_s_1_2_2(or_822_cse, or_361_cse, fsm_output[6]);
  assign mux_623_cse = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), fsm_output[7]);
  assign mux_624_cse = MUX_s_1_2_2(mux_623_cse, or_361_cse, fsm_output[6]);
  assign or_tmp_611 = (fsm_output[1]) | (fsm_output[0]) | (fsm_output[2]) | (~ (fsm_output[4]));
  assign nand_163_cse = ~(reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1 & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1);
  assign or_dcpl_770 = (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2)
      | reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0;
  assign or_1420_cse = reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1 | reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  assign or_dcpl_774 = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 | reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0;
  assign or_1431_cse = (~ reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1) | reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  assign or_1435_cse = reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1 | (~ reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1);
  assign or_dcpl_791 = ~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 &
      reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0);
  assign or_dcpl_794 = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 | (~
      reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0);
  assign and_dcpl_148 = (fsm_output[7:6]==2'b11);
  assign or_tmp_682 = (fsm_output[5:4]!=2'b01);
  assign or_dcpl_959 = ~((fsm_output[8]) & (fsm_output[4]));
  assign or_dcpl_961 = or_dcpl_959 | (~ (fsm_output[2])) | nand_197_cse;
  assign and_dcpl_181 = (~ (fsm_output[5])) & (fsm_output[3]);
  assign and_dcpl_182 = and_dcpl_181 & and_dcpl_148;
  assign and_dcpl_185 = and_dcpl_61 & (~ (fsm_output[2]));
  assign and_dcpl_186 = and_dcpl_185 & nor_777_cse;
  assign and_dcpl_187 = and_dcpl_186 & and_dcpl_182;
  assign and_dcpl_189 = (fsm_output[5]) & (~ (fsm_output[3]));
  assign and_dcpl_190 = and_dcpl_189 & and_dcpl_45;
  assign and_dcpl_191 = and_dcpl_61 & (fsm_output[2]);
  assign and_dcpl_192 = and_dcpl_191 & nor_777_cse;
  assign and_dcpl_193 = and_dcpl_192 & and_dcpl_190;
  assign and_dcpl_194 = (fsm_output[5]) & (fsm_output[3]);
  assign and_dcpl_197 = and_dcpl_186 & and_dcpl_194 & (~ (z_out_5[2])) & and_dcpl_45;
  assign and_dcpl_198 = ~((fsm_output[5]) | (fsm_output[3]));
  assign and_dcpl_199 = and_dcpl_198 & and_dcpl_45;
  assign and_dcpl_200 = (fsm_output[1:0]==2'b01);
  assign and_dcpl_201 = (~ (fsm_output[8])) & (fsm_output[4]);
  assign and_dcpl_202 = and_dcpl_201 & (fsm_output[2]);
  assign and_dcpl_203 = and_dcpl_202 & and_dcpl_200;
  assign and_dcpl_204 = and_dcpl_203 & and_dcpl_199;
  assign or_dcpl_980 = or_dcpl_512 | or_dcpl_4;
  assign or_dcpl_983 = or_76_cse | or_dcpl_96;
  assign or_dcpl_985 = or_dcpl_508 | or_dcpl_4;
  assign or_dcpl_987 = or_130_cse | or_dcpl_96;
  assign or_dcpl_988 = or_130_cse | or_dcpl_4;
  assign or_dcpl_989 = or_dcpl_508 | or_dcpl_96;
  assign or_dcpl_990 = or_76_cse | or_dcpl_4;
  assign or_dcpl_991 = or_dcpl_512 | or_dcpl_96;
  assign or_dcpl_993 = or_dcpl_512 | or_dcpl_584;
  assign or_dcpl_995 = or_76_cse | or_dcpl_54;
  assign or_dcpl_996 = or_dcpl_508 | or_dcpl_584;
  assign or_dcpl_997 = or_130_cse | or_dcpl_54;
  assign or_dcpl_998 = or_130_cse | or_dcpl_584;
  assign or_dcpl_999 = or_dcpl_508 | or_dcpl_54;
  assign or_dcpl_1000 = or_dcpl_512 | or_dcpl_54;
  assign and_dcpl_205 = and_dcpl_201 & (~ (fsm_output[2]));
  assign and_dcpl_206 = and_dcpl_205 & and_dcpl_200;
  assign and_dcpl_207 = and_dcpl_206 & and_dcpl_199;
  assign or_dcpl_1001 = ~(reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1);
  assign or_dcpl_1002 = or_130_cse | or_dcpl_1001;
  assign or_dcpl_1003 = reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 | reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  assign or_dcpl_1004 = or_dcpl_508 | or_dcpl_1003;
  assign or_dcpl_1005 = (~ reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0) | reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  assign or_dcpl_1006 = or_130_cse | or_dcpl_1005;
  assign or_dcpl_1007 = reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 | (~ reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1);
  assign or_dcpl_1008 = or_dcpl_508 | or_dcpl_1007;
  assign or_dcpl_1009 = or_130_cse | or_dcpl_1007;
  assign or_dcpl_1010 = or_dcpl_508 | or_dcpl_1005;
  assign or_dcpl_1011 = or_130_cse | or_dcpl_1003;
  assign or_dcpl_1012 = or_dcpl_508 | or_dcpl_1001;
  assign or_dcpl_1013 = or_76_cse | or_dcpl_1001;
  assign or_dcpl_1014 = or_dcpl_512 | or_dcpl_1003;
  assign or_dcpl_1015 = or_76_cse | or_dcpl_1005;
  assign or_dcpl_1016 = or_dcpl_512 | or_dcpl_1007;
  assign or_dcpl_1017 = or_76_cse | or_dcpl_1007;
  assign or_dcpl_1018 = or_dcpl_512 | or_dcpl_1005;
  assign or_dcpl_1019 = or_dcpl_512 | or_dcpl_1001;
  assign and_dcpl_209 = and_dcpl_198 & nor_973_cse;
  assign and_dcpl_211 = (fsm_output[1:0]==2'b10);
  assign and_dcpl_212 = and_dcpl_205 & and_dcpl_211;
  assign and_dcpl_213 = and_dcpl_212 & and_dcpl_199;
  assign nor_tmp_261 = ((~((fsm_output[2]) | (~ (fsm_output[6])))) | (fsm_output[4]))
      & (fsm_output[7]);
  assign and_dcpl_215 = and_dcpl_202 & and_dcpl_211;
  assign and_dcpl_216 = and_dcpl_215 & and_dcpl_199;
  assign mux_tmp_787 = MUX_s_1_2_2((~ (fsm_output[1])), (fsm_output[1]), fsm_output[0]);
  assign mux_tmp_788 = MUX_s_1_2_2(nand_197_cse, mux_tmp_787, fsm_output[3]);
  assign and_dcpl_220 = (~ mux_tmp_788) & and_dcpl_61 & (~((fsm_output[2]) | (fsm_output[5])))
      & and_dcpl_148;
  assign and_dcpl_221 = and_dcpl_198 & and_dcpl_148;
  assign and_dcpl_222 = and_dcpl_192 & and_dcpl_221;
  assign or_dcpl_1020 = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 | (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd);
  assign or_dcpl_1021 = or_dcpl_1020 | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign or_dcpl_1022 = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd;
  assign or_dcpl_1023 = or_dcpl_1022 | (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign or_dcpl_1024 = or_dcpl_1020 | (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign and_dcpl_226 = ~((fsm_output[8]) | (fsm_output[2]));
  assign or_tmp_704 = (fsm_output[1]) | (fsm_output[4]);
  assign nand_253_cse = ~((fsm_output[7:6]==2'b11));
  assign or_tmp_708 = (fsm_output[3]) | nand_253_cse;
  assign and_dcpl_231 = (fsm_output[3]) & (fsm_output[6]);
  assign or_dcpl_1025 = or_76_cse | or_dcpl_584;
  assign and_dcpl_237 = and_dcpl_181 & and_dcpl_45;
  assign and_dcpl_239 = and_dcpl_191 & and_1474_cse;
  assign and_dcpl_240 = and_dcpl_239 & and_dcpl_237;
  assign or_dcpl_1026 = ~(reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd);
  assign or_dcpl_1027 = (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1) | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd;
  assign or_dcpl_1028 = or_dcpl_1027 | or_dcpl_1026;
  assign or_dcpl_1029 = reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 | reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd;
  assign or_dcpl_1030 = or_dcpl_1020 | or_dcpl_1029;
  assign or_dcpl_1031 = or_dcpl_1022 | or_dcpl_1026;
  assign or_dcpl_1032 = ~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd);
  assign or_dcpl_1033 = or_dcpl_1032 | or_dcpl_1029;
  assign or_dcpl_1034 = (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1) |
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd;
  assign or_dcpl_1035 = or_dcpl_1027 | or_dcpl_1034;
  assign or_dcpl_1036 = reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 | (~
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd);
  assign or_dcpl_1037 = or_dcpl_1020 | or_dcpl_1036;
  assign or_dcpl_1038 = or_dcpl_1022 | or_dcpl_1034;
  assign or_dcpl_1039 = or_dcpl_1032 | or_dcpl_1036;
  assign or_dcpl_1040 = or_dcpl_1027 | or_dcpl_1036;
  assign or_dcpl_1041 = or_dcpl_1020 | or_dcpl_1034;
  assign or_dcpl_1042 = or_dcpl_1022 | or_dcpl_1036;
  assign or_dcpl_1043 = or_dcpl_1032 | or_dcpl_1034;
  assign or_dcpl_1044 = or_dcpl_1027 | or_dcpl_1029;
  assign or_dcpl_1045 = or_dcpl_1020 | or_dcpl_1026;
  assign or_dcpl_1046 = or_dcpl_1032 | or_dcpl_1026;
  assign and_dcpl_241 = and_dcpl_185 & and_1474_cse;
  assign and_dcpl_242 = and_dcpl_241 & and_dcpl_209;
  assign and_dcpl_243 = (fsm_output[3]) & (~ (fsm_output[6]));
  assign and_dcpl_248 = and_dcpl_205 & and_dcpl_200 & (fsm_output[5]) & and_dcpl_243
      & (~ (fsm_output[7])) & (~((RMS_NORM_LOOP_2_2_i_4_0_sva_1[4]) & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1));
  assign and_dcpl_252 = (fsm_output[8]) & (~ (fsm_output[4]));
  assign and_dcpl_255 = and_dcpl_252 & (~ (fsm_output[2])) & nor_777_cse & and_dcpl_198
      & and_dcpl_57;
  assign and_dcpl_256 = and_dcpl_181 & and_dcpl_57;
  assign and_dcpl_257 = and_dcpl_239 & and_dcpl_256;
  assign and_dcpl_258 = (~ (fsm_output[8])) & (fsm_output[6]);
  assign and_dcpl_259 = and_dcpl_258 & (~ (fsm_output[7]));
  assign or_tmp_728 = and_1559_cse | (fsm_output[4]);
  assign mux_817_nl = MUX_s_1_2_2((~ (fsm_output[4])), or_tmp_728, fsm_output[5]);
  assign mux_819_nl = MUX_s_1_2_2(mux_tmp_91, mux_817_nl, fsm_output[3]);
  assign and_dcpl_260 = (~ mux_819_nl) & and_dcpl_259;
  assign mux_tmp_824 = MUX_s_1_2_2(mux_tmp_121, or_2456_cse, fsm_output[4]);
  assign nand_257_nl = ~((fsm_output[6]) & (fsm_output[8]));
  assign mux_827_nl = MUX_s_1_2_2(nand_257_nl, or_tmp_464, fsm_output[4]);
  assign mux_828_nl = MUX_s_1_2_2(mux_827_nl, or_2742_cse, fsm_output[0]);
  assign mux_829_nl = MUX_s_1_2_2(mux_828_nl, mux_tmp_824, fsm_output[5]);
  assign or_1090_nl = (fsm_output[3:2]!=2'b00);
  assign mux_830_nl = MUX_s_1_2_2(mux_829_nl, mux_2032_cse, or_1090_nl);
  assign mux_822_nl = MUX_s_1_2_2(or_2742_cse, mux_2024_cse, fsm_output[0]);
  assign mux_823_nl = MUX_s_1_2_2(mux_822_nl, or_2736_cse, fsm_output[5]);
  assign mux_826_nl = MUX_s_1_2_2(mux_2032_cse, mux_823_nl, and_1773_cse);
  assign mux_831_nl = MUX_s_1_2_2(mux_830_nl, mux_826_nl, fsm_output[1]);
  assign or_dcpl_1048 = mux_831_nl | (fsm_output[7]);
  assign and_dcpl_261 = and_dcpl_181 & nor_973_cse;
  assign and_dcpl_263 = nor_tmp_99 & (fsm_output[2]);
  assign and_dcpl_264 = and_dcpl_263 & and_1474_cse;
  assign and_dcpl_265 = and_dcpl_264 & and_dcpl_261;
  assign or_dcpl_1050 = ~((fsm_output[4]) & (fsm_output[2]));
  assign and_dcpl_268 = (or_dcpl_1050 | (~((fsm_output[1]) & (fsm_output[3])))) &
      (fsm_output[8]) & (fsm_output[5]) & nor_973_cse;
  assign and_dcpl_270 = and_dcpl_1 & nor_973_cse;
  assign mux_tmp_834 = MUX_s_1_2_2(or_tmp_11, or_270_cse, fsm_output[1]);
  assign mux_833_nl = MUX_s_1_2_2(mux_tmp_87, or_270_cse, fsm_output[1]);
  assign mux_835_nl = MUX_s_1_2_2(mux_tmp_834, mux_833_nl, fsm_output[0]);
  assign mux_tmp_836 = MUX_s_1_2_2(mux_835_nl, (fsm_output[4]), fsm_output[3]);
  assign and_dcpl_272 = (~ (fsm_output[8])) & (fsm_output[2]);
  assign and_dcpl_275 = and_dcpl_194 & nor_973_cse;
  assign and_dcpl_276 = and_dcpl_212 & and_dcpl_275;
  assign or_3137_cse = and_1474_cse | (fsm_output[2]);
  assign nor_tmp_282 = or_3137_cse & (fsm_output[4]);
  assign and_1498_nl = (fsm_output[3]) & (fsm_output[5]) & nor_tmp_282;
  assign nor_897_nl = ~((fsm_output[5:3]!=3'b000));
  assign mux_837_nl = MUX_s_1_2_2(and_1498_nl, nor_897_nl, fsm_output[6]);
  assign and_dcpl_278 = mux_837_nl & and_dcpl_26;
  assign and_dcpl_279 = (fsm_output[5:4]==2'b01);
  assign or_tmp_742 = (fsm_output[7]) | (fsm_output[5]) | (fsm_output[8]);
  assign mux_tmp_839 = MUX_s_1_2_2(or_tmp_742, or_1767_cse, fsm_output[4]);
  assign or_1795_cse = (fsm_output[7]) | (~ (fsm_output[5])) | (fsm_output[8]);
  assign mux_tmp_841 = MUX_s_1_2_2(or_tmp_742, or_1795_cse, fsm_output[4]);
  assign nor_tmp_285 = or_3185_cse & (fsm_output[4]);
  assign and_dcpl_289 = and_dcpl_202 & nor_777_cse;
  assign and_dcpl_290 = and_dcpl_289 & and_dcpl_209;
  assign and_dcpl_291 = and_dcpl_189 & and_dcpl_148;
  assign and_dcpl_292 = and_dcpl_186 & and_dcpl_291;
  assign and_dcpl_293 = and_dcpl_194 & and_dcpl_45;
  assign and_dcpl_294 = and_dcpl_239 & and_dcpl_293;
  assign and_dcpl_295 = (fsm_output[8:7]==2'b01);
  assign or_tmp_755 = (fsm_output[5:1]!=5'b00000);
  assign and_dcpl_298 = (~ (fsm_output[8])) & (fsm_output[5]) & and_dcpl_148;
  assign and_dcpl_302 = and_dcpl_194 & and_dcpl_148;
  assign or_tmp_757 = nor_717_cse | (~ (fsm_output[4])) | (fsm_output[8]);
  assign or_tmp_762 = and_1572_cse | (fsm_output[4]);
  assign and_337_nl = (fsm_output[5]) & or_tmp_762;
  assign mux_tmp_857 = MUX_s_1_2_2(and_1762_cse, and_337_nl, fsm_output[3]);
  assign mux_858_nl = MUX_s_1_2_2(mux_tmp_857, (~ or_tmp_755), fsm_output[6]);
  assign and_dcpl_304 = mux_858_nl & and_dcpl_295;
  assign nor_tmp_289 = or_1908_cse & (fsm_output[4]);
  assign and_dcpl_306 = and_dcpl_264 & and_dcpl_275;
  assign and_dcpl_307 = ~((fsm_output[8]) | (fsm_output[6]));
  assign and_dcpl_308 = and_dcpl_307 & (~ (fsm_output[7]));
  assign nor_tmp_291 = or_1732_cse & (fsm_output[2]) & (fsm_output[4]);
  assign or_tmp_767 = and_1637_cse | (fsm_output[4]);
  assign and_344_nl = (fsm_output[5]) & or_tmp_728;
  assign mux_866_nl = MUX_s_1_2_2(and_1762_cse, and_344_nl, fsm_output[3]);
  assign nand_262_nl = ~((fsm_output[6]) & mux_866_nl);
  assign or_1827_nl = (fsm_output[5]) | or_tmp_767;
  assign mux_865_nl = MUX_s_1_2_2(or_2699_cse, or_1827_nl, fsm_output[3]);
  assign or_3142_nl = (fsm_output[6]) | mux_865_nl;
  assign mux_867_nl = MUX_s_1_2_2(nand_262_nl, or_3142_nl, fsm_output[7]);
  assign and_dcpl_310 = ~(mux_867_nl | (fsm_output[8]));
  assign and_dcpl_312 = and_dcpl_185 & and_dcpl_200;
  assign and_dcpl_313 = and_dcpl_312 & and_dcpl_190;
  assign and_dcpl_315 = and_dcpl_191 & and_dcpl_200;
  assign and_dcpl_316 = and_dcpl_315 & and_dcpl_221;
  assign and_dcpl_318 = and_dcpl_202 & and_1474_cse & and_dcpl_199;
  assign and_dcpl_319 = and_dcpl & (fsm_output[7]);
  assign and_dcpl_321 = and_1474_cse & (~ (fsm_output[5]));
  assign and_dcpl_322 = and_dcpl_202 & and_dcpl_321;
  assign and_dcpl_327 = and_dcpl_205 & and_1474_cse;
  assign and_dcpl_328 = and_dcpl_327 & and_dcpl_237;
  assign or_1835_cse = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[5]);
  assign and_dcpl_334 = ~((reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1!=2'b00));
  assign and_dcpl_335 = and_dcpl_334 & (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  assign and_dcpl_336 = nor_973_cse & (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd);
  assign and_dcpl_338 = (fsm_output[0]) & (~ (fsm_output[5]));
  assign and_dcpl_339 = and_dcpl_338 & (~ (fsm_output[3]));
  assign and_dcpl_341 = and_dcpl_61 & nor_717_cse;
  assign and_dcpl_342 = and_dcpl_341 & and_dcpl_339;
  assign nor_tmp_307 = (fsm_output[5]) & (fsm_output[8]);
  assign and_dcpl_344 = and_dcpl_206 & and_dcpl_275;
  assign and_dcpl_346 = and_dcpl_201 & and_dcpl_211 & and_dcpl_199;
  assign nand_263_cse = ~((fsm_output[0]) & (fsm_output[1]) & (fsm_output[4]));
  assign or_tmp_798 = (fsm_output[5]) | nand_263_cse;
  assign mux_903_nl = MUX_s_1_2_2(or_1867_cse, or_tmp_704, fsm_output[0]);
  assign nand_44_nl = ~((fsm_output[5]) & (~ mux_903_nl));
  assign mux_904_nl = MUX_s_1_2_2(nand_44_nl, or_tmp_798, fsm_output[3]);
  assign and_dcpl_348 = (~ mux_904_nl) & and_dcpl_272 & and_dcpl_45;
  assign and_dcpl_349 = and_dcpl_312 & and_dcpl_293;
  assign and_dcpl_350 = and_dcpl_185 & and_dcpl_211;
  assign and_dcpl_351 = and_dcpl_350 & and_dcpl_221;
  assign and_dcpl_352 = and_dcpl_241 & and_dcpl_182;
  assign and_dcpl_353 = ~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2]) | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]));
  assign and_dcpl_354 = and_dcpl_353 & (~ reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  assign and_dcpl_355 = and_dcpl_148 & (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[1]));
  assign and_dcpl_357 = (fsm_output[0]) & (fsm_output[5]);
  assign and_dcpl_360 = and_dcpl_201 & and_1559_cse & and_dcpl_357 & (~ (fsm_output[3]));
  assign or_dcpl_1063 = or_dcpl_774 | or_1420_cse;
  assign and_dcpl_362 = and_dcpl_205 & nor_777_cse;
  assign and_dcpl_363 = and_dcpl_362 & and_dcpl_275;
  assign and_dcpl_364 = (fsm_output[4]) & (~ (fsm_output[2]));
  assign and_dcpl_374 = and_dcpl_201 & nor_717_cse & and_dcpl_339 & and_dcpl_45 &
      (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1) & (~(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1));
  assign or_tmp_805 = (~((fsm_output[7:6]!=2'b01))) | (fsm_output[8]);
  assign mux_tmp_906 = MUX_s_1_2_2(or_362_cse, or_361_cse, fsm_output[6]);
  assign or_tmp_808 = (fsm_output[8:6]!=3'b000);
  assign mux_tmp_908 = MUX_s_1_2_2(or_1197_cse, or_tmp_808, fsm_output[4]);
  assign mux_tmp_910 = MUX_s_1_2_2(mux_tmp_604, or_tmp_808, fsm_output[4]);
  assign or_tmp_812 = (fsm_output[8:6]!=3'b010);
  assign mux_tmp_915 = MUX_s_1_2_2(mux_tmp_906, or_tmp_812, fsm_output[4]);
  assign or_tmp_813 = (fsm_output[6]) | ((fsm_output[8:7]==2'b11));
  assign mux_tmp_916 = MUX_s_1_2_2(or_822_cse, (fsm_output[8]), fsm_output[6]);
  assign mux_tmp_919 = MUX_s_1_2_2(or_822_cse, or_362_cse, fsm_output[6]);
  assign or_tmp_814 = (fsm_output[6]) | mux_623_cse;
  assign mux_tmp_922 = MUX_s_1_2_2(mux_tmp_919, or_tmp_814, fsm_output[4]);
  assign mux_tmp_927 = MUX_s_1_2_2(mux_tmp_906, or_tmp_805, fsm_output[4]);
  assign mux_tmp_936 = MUX_s_1_2_2((fsm_output[7]), or_362_cse, fsm_output[6]);
  assign mux_tmp_937 = MUX_s_1_2_2(mux_tmp_936, or_tmp_814, fsm_output[4]);
  assign and_dcpl_376 = and_dcpl_191 & and_dcpl_211;
  assign and_dcpl_377 = and_dcpl_376 & and_dcpl_293;
  assign or_3149_nl = (fsm_output[6]) | (~ (fsm_output[2])) | (fsm_output[4]);
  assign or_3150_nl = (~ (fsm_output[6])) | (fsm_output[2]) | (~ (fsm_output[4]));
  assign mux_953_nl = MUX_s_1_2_2(or_3149_nl, or_3150_nl, fsm_output[7]);
  assign and_dcpl_381 = ~(mux_953_nl | (fsm_output[8]));
  assign and_dcpl_382 = and_dcpl_381 & and_dcpl_200 & and_dcpl_198;
  assign or_tmp_833 = (~ (fsm_output[2])) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign nor_923_nl = ~((~((fsm_output[2]) | (~ (fsm_output[4])))) | (fsm_output[8]));
  assign nand_264_nl = ~(or_dcpl_1050 & (fsm_output[8]));
  assign mux_tmp_960 = MUX_s_1_2_2(nor_923_nl, nand_264_nl, fsm_output[1]);
  assign mux_tmp_967 = MUX_s_1_2_2(or_tmp_48, or_133_cse, fsm_output[2]);
  assign or_1910_nl = (fsm_output[2]) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_tmp_968 = MUX_s_1_2_2(or_1910_nl, mux_tmp_967, fsm_output[1]);
  assign and_dcpl_383 = (fsm_output[2:1]==2'b10);
  assign or_1912_nl = (fsm_output[6]) | (~ (fsm_output[0]));
  assign or_3073_nl = (~ (fsm_output[6])) | (fsm_output[0]);
  assign mux_tmp_975 = MUX_s_1_2_2(or_1912_nl, or_3073_nl, fsm_output[7]);
  assign and_dcpl_385 = (~ mux_tmp_975) & and_dcpl_201;
  assign and_dcpl_386 = and_dcpl_385 & and_dcpl_383 & and_dcpl_189;
  assign and_dcpl_388 = and_dcpl_1 & (fsm_output[7]);
  assign or_tmp_861 = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[2]) | (fsm_output[4]);
  assign and_dcpl_390 = and_dcpl_226 & and_dcpl_45;
  assign or_tmp_878 = ~((fsm_output[0]) & (fsm_output[1]) & (fsm_output[4]) & (~
      (fsm_output[8])));
  assign and_dcpl_410 = and_dcpl_376 & and_dcpl_237;
  assign and_dcpl_413 = (fsm_output[8:6]==3'b100);
  assign nor_tmp_329 = (fsm_output[0]) & (fsm_output[1]) & (fsm_output[2]) & (fsm_output[4]);
  assign mux_1026_nl = MUX_s_1_2_2((~ nor_tmp_285), nor_tmp_329, fsm_output[5]);
  assign mux_tmp_1027 = MUX_s_1_2_2((~ (fsm_output[5])), mux_1026_nl, fsm_output[3]);
  assign and_dcpl_414 = (~ mux_tmp_1027) & and_dcpl_413;
  assign and_dcpl_415 = and_dcpl_312 & and_dcpl_209;
  assign or_1976_nl = (fsm_output[5]) | (fsm_output[2]) | (~ (fsm_output[4]));
  assign or_1974_nl = (fsm_output[5]) | (~ (fsm_output[1])) | (~ (fsm_output[2]))
      | (fsm_output[4]);
  assign mux_1028_nl = MUX_s_1_2_2(or_1976_nl, or_1974_nl, fsm_output[3]);
  assign or_tmp_913 = (fsm_output[6]) | mux_1028_nl;
  assign or_tmp_914 = (fsm_output[7:5]!=3'b010);
  assign and_dcpl_417 = nor_973_cse & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd;
  assign and_dcpl_420 = and_dcpl & (~ (fsm_output[7]));
  assign and_dcpl_421 = and_dcpl_200 & (~ (fsm_output[5]));
  assign and_dcpl_422 = and_dcpl_421 & and_dcpl_420;
  assign or_dcpl_1067 = or_619_cse | or_750_cse;
  assign and_dcpl_425 = and_dcpl_189 & nor_973_cse;
  assign or_tmp_922 = (fsm_output[4]) | (~ (fsm_output[7]));
  assign or_tmp_923 = (~ (fsm_output[4])) | (fsm_output[7]);
  assign mux_tmp_1044 = MUX_s_1_2_2((~ or_tmp_923), or_tmp_922, fsm_output[5]);
  assign or_tmp_930 = (fsm_output[5]) | (fsm_output[4]) | (~ (fsm_output[7]));
  assign mux_tmp_1051 = MUX_s_1_2_2(or_tmp_922, or_tmp_923, fsm_output[5]);
  assign mux_tmp_1052 = MUX_s_1_2_2((~ (fsm_output[7])), or_tmp_923, fsm_output[5]);
  assign or_tmp_931 = (fsm_output[5]) | (~ (fsm_output[7]));
  assign or_dcpl_1068 = or_dcpl_1022 | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign and_dcpl_432 = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1==2'b01);
  assign and_dcpl_433 = and_dcpl_432 & (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  assign or_dcpl_1070 = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1]);
  assign or_dcpl_1071 = or_dcpl_1070 | or_790_cse;
  assign and_dcpl_438 = and_dcpl_203 & and_dcpl_425;
  assign and_dcpl_439 = and_dcpl_312 & and_dcpl_256;
  assign or_tmp_938 = (fsm_output[5]) | (fsm_output[3]) | (~ (fsm_output[7]));
  assign not_tmp_549 = ~((fsm_output[5]) & (fsm_output[3]) & (fsm_output[7]));
  assign and_dcpl_442 = and_dcpl_350 & and_dcpl_293;
  assign and_dcpl_448 = and_dcpl_289 & and_dcpl_291;
  assign and_dcpl_449 = nor_tmp_99 & (~ (fsm_output[2]));
  assign and_dcpl_452 = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1==2'b10);
  assign and_dcpl_453 = and_dcpl_452 & (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  assign or_dcpl_1073 = nand_143_cse | or_750_cse;
  assign and_dcpl_458 = and_dcpl_353 & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1;
  assign or_dcpl_1076 = or_dcpl_770 | or_1435_cse;
  assign and_dcpl_461 = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1==2'b11);
  assign and_dcpl_462 = and_dcpl_461 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  assign or_dcpl_1077 = ~((reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0])
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  assign or_dcpl_1079 = or_806_cse | or_dcpl_1077;
  assign and_dcpl_467 = (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2]) & (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]);
  assign and_dcpl_468 = and_dcpl_467 & (~ reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  assign or_dcpl_1081 = or_dcpl_774 | or_1431_cse;
  assign and_dcpl_471 = and_dcpl_452 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  assign or_dcpl_1083 = nand_143_cse | or_753_cse;
  assign and_dcpl_477 = and_dcpl_385 & nor_717_cse & and_dcpl_194;
  assign and_dcpl_478 = and_dcpl_1 & (~ (fsm_output[3]));
  assign or_tmp_992 = nor_777_cse | (~ (fsm_output[2])) | (fsm_output[4]);
  assign mux_tmp_1113 = MUX_s_1_2_2(or_dcpl_1050, or_tmp_11, fsm_output[1]);
  assign or_tmp_993 = (fsm_output[6]) | (fsm_output[0]) | (~ (fsm_output[1])) | (fsm_output[2])
      | (fsm_output[4]);
  assign and_dcpl_480 = and_dcpl_334 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  assign or_dcpl_1084 = or_dcpl_1070 | or_753_cse;
  assign and_dcpl_486 = and_dcpl_461 & (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2);
  assign or_dcpl_1085 = nand_143_cse | or_790_cse;
  assign or_dcpl_1086 = or_806_cse | or_790_cse;
  assign or_dcpl_1087 = or_619_cse | or_753_cse;
  assign or_dcpl_1088 = or_806_cse | or_753_cse;
  assign or_dcpl_1089 = or_619_cse | or_790_cse;
  assign mux_tmp_1120 = MUX_s_1_2_2(or_2456_cse, or_tmp_464, fsm_output[7]);
  assign mux_1122_cse = MUX_s_1_2_2(or_1197_cse, mux_tmp_1120, fsm_output[4]);
  assign mux_1125_cse = MUX_s_1_2_2(or_1197_cse, mux_502_cse, fsm_output[4]);
  assign and_dcpl_511 = (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2]) & (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]));
  assign and_dcpl_512 = and_dcpl_511 & (~ reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  assign and_dcpl_513 = and_dcpl_148 & (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[1]);
  assign or_dcpl_1090 = or_806_cse | or_750_cse;
  assign mux_1148_nl = MUX_s_1_2_2(nand_197_cse, or_2792_cse, fsm_output[3]);
  assign mux_1149_nl = MUX_s_1_2_2(mux_tmp_788, mux_1148_nl, z_out_5[2]);
  assign and_dcpl_524 = (~(mux_1149_nl | (fsm_output[8]))) & nor_992_cse & (~ (fsm_output[5]))
      & and_dcpl_148;
  assign nor_354_cse = ~((fsm_output[3]) | (~ (fsm_output[1])));
  assign nor_355_cse = ~((fsm_output[1:0]!=2'b10) | (~ (z_out_5[2])));
  assign mux_1158_nl = MUX_s_1_2_2(or_1197_cse, or_1984_cse, fsm_output[1]);
  assign mux_1157_nl = MUX_s_1_2_2(or_1984_cse, mux_tmp_1120, fsm_output[1]);
  assign mux_1159_nl = MUX_s_1_2_2(mux_1158_nl, mux_1157_nl, fsm_output[0]);
  assign mux_1156_nl = MUX_s_1_2_2(mux_tmp_1120, or_1197_cse, nor_355_cse);
  assign mux_1160_nl = MUX_s_1_2_2(mux_1159_nl, mux_1156_nl, fsm_output[3]);
  assign mux_1161_nl = MUX_s_1_2_2(mux_1160_nl, mux_tmp_1120, fsm_output[2]);
  assign mux_1154_nl = MUX_s_1_2_2(mux_tmp_1120, mux_502_cse, nor_354_cse);
  assign mux_1152_nl = MUX_s_1_2_2(mux_502_cse, mux_tmp_1120, and_1474_cse);
  assign mux_1153_nl = MUX_s_1_2_2(mux_1152_nl, or_tmp_507, fsm_output[3]);
  assign mux_1155_nl = MUX_s_1_2_2(mux_1154_nl, mux_1153_nl, fsm_output[2]);
  assign mux_1162_nl = MUX_s_1_2_2(mux_1161_nl, mux_1155_nl, fsm_output[4]);
  assign mux_tmp_1163 = MUX_s_1_2_2(mux_1162_nl, or_tmp_507, fsm_output[5]);
  assign and_dcpl_525 = and_dcpl_511 & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1;
  assign and_dcpl_528 = and_dcpl_432 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2;
  assign or_dcpl_1091 = or_619_cse | or_dcpl_1077;
  assign or_dcpl_1092 = or_dcpl_1070 | or_dcpl_1077;
  assign mux_tmp_1178 = MUX_s_1_2_2(or_2455_cse, or_tmp_464, fsm_output[7]);
  assign mux_tmp_1179 = MUX_s_1_2_2(mux_tmp_1178, or_tmp_507, fsm_output[4]);
  assign mux_tmp_1183 = MUX_s_1_2_2((fsm_output[6]), or_tmp_464, fsm_output[7]);
  assign mux_tmp_1185 = MUX_s_1_2_2(or_1984_cse, mux_tmp_1183, fsm_output[4]);
  assign mux_tmp_1187 = MUX_s_1_2_2((fsm_output[6]), (fsm_output[8]), fsm_output[7]);
  assign or_tmp_1035 = and_1474_cse | (fsm_output[3]) | (fsm_output[8]);
  assign and_dcpl_539 = and_dcpl_467 & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1;
  assign or_tmp_1051 = (~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[8]));
  assign mux_tmp_1218 = MUX_s_1_2_2(or_362_cse, or_822_cse, fsm_output[5]);
  assign mux_tmp_1219 = MUX_s_1_2_2((fsm_output[8]), or_822_cse, fsm_output[5]);
  assign mux_tmp_1229 = MUX_s_1_2_2(or_361_cse, or_822_cse, fsm_output[5]);
  assign mux_tmp_1237 = MUX_s_1_2_2(nand_253_cse, or_1984_cse, fsm_output[8]);
  assign mux_tmp_1238 = MUX_s_1_2_2(mux_tmp_1237, or_1197_cse, fsm_output[5]);
  assign or_tmp_1066 = (fsm_output[8]) | nand_253_cse;
  assign mux_tmp_1240 = MUX_s_1_2_2(or_tmp_1066, or_1197_cse, fsm_output[5]);
  assign mux_tmp_1245 = MUX_s_1_2_2(or_tmp_808, or_1197_cse, fsm_output[5]);
  assign mux_1249_nl = MUX_s_1_2_2(mux_792_cse, or_1984_cse, fsm_output[8]);
  assign mux_tmp_1250 = MUX_s_1_2_2(or_tmp_1066, mux_1249_nl, fsm_output[5]);
  assign and_dcpl_548 = and_dcpl_362 & and_dcpl_302;
  assign and_dcpl_549 = ~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd |
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[1]));
  assign and_dcpl_550 = and_dcpl_549 & (~ (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]));
  assign and_dcpl_551 = nor_973_cse & (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1);
  assign and_dcpl_552 = and_dcpl_551 & and_dcpl_550;
  assign and_dcpl_553 = and_dcpl_338 & (fsm_output[3]);
  assign and_dcpl_554 = (fsm_output[2:1]==2'b01);
  assign and_dcpl_557 = nor_tmp_99 & and_dcpl_554 & and_dcpl_553 & and_dcpl_552;
  assign mux_tmp_1281 = MUX_s_1_2_2(or_255_cse, or_270_cse, fsm_output[1]);
  assign and_dcpl_564 = and_dcpl_198 & (~ (fsm_output[6]));
  assign and_dcpl_576 = (fsm_output[3]) & (~ (fsm_output[7]));
  assign and_dcpl_577 = ~((fsm_output[1]) | (fsm_output[5]));
  assign mux_1309_cse = MUX_s_1_2_2(or_dcpl_959, or_133_cse, fsm_output[6]);
  assign and_dcpl_581 = and_dcpl_1 & and_dcpl_45;
  assign or_tmp_1128 = (~ (fsm_output[1])) | (~ (fsm_output[2])) | (fsm_output[4]);
  assign and_dcpl_583 = and_dcpl_327 & and_dcpl_199;
  assign or_2235_nl = (fsm_output[5]) | or_tmp_762;
  assign mux_1311_nl = MUX_s_1_2_2(or_2699_cse, or_2235_nl, fsm_output[3]);
  assign or_tmp_1132 = (fsm_output[6]) | mux_1311_nl;
  assign and_443_nl = (fsm_output[5]) & nor_tmp_291;
  assign mux_1312_nl = MUX_s_1_2_2(and_443_nl, and_1762_cse, fsm_output[3]);
  assign nor_930_nl = ~((fsm_output[6]) | mux_1312_nl);
  assign mux_1313_nl = MUX_s_1_2_2(nor_930_nl, or_tmp_1132, fsm_output[7]);
  assign or_dcpl_1104 = mux_1313_nl | (fsm_output[8]);
  assign and_dcpl_585 = and_dcpl_57 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd;
  assign and_dcpl_586 = and_dcpl_585 & and_dcpl_486;
  assign and_dcpl_587 = and_dcpl_61 & and_dcpl_554;
  assign and_dcpl_588 = and_dcpl_587 & and_dcpl_553;
  assign and_dcpl_591 = and_dcpl_57 & (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd);
  assign and_dcpl_592 = and_dcpl_591 & and_dcpl_480;
  assign and_dcpl_595 = and_dcpl_585 & and_dcpl_471;
  assign and_dcpl_598 = and_dcpl_591 & and_dcpl_433;
  assign and_dcpl_601 = and_dcpl_585 & and_dcpl_453;
  assign and_dcpl_604 = and_dcpl_591 & and_dcpl_528;
  assign and_dcpl_607 = and_dcpl_585 & and_dcpl_528;
  assign and_dcpl_610 = and_dcpl_591 & and_dcpl_453;
  assign and_dcpl_613 = and_dcpl_585 & and_dcpl_433;
  assign and_dcpl_616 = and_dcpl_591 & and_dcpl_471;
  assign mux_1396_nl = MUX_s_1_2_2(or_2249_cse, or_1983_cse, fsm_output[2]);
  assign and_1616_nl = (fsm_output[3]) & (fsm_output[0]) & (fsm_output[1]);
  assign mux_1398_nl = MUX_s_1_2_2(mux_806_cse, mux_1396_nl, and_1616_nl);
  assign mux_1399_nl = MUX_s_1_2_2(mux_1398_nl, or_1983_cse, fsm_output[5]);
  assign or_2296_nl = (~(and_1637_cse | (fsm_output[6]))) | (fsm_output[7]);
  assign mux_1394_nl = MUX_s_1_2_2(or_2296_nl, (fsm_output[7]), fsm_output[3]);
  assign mux_1395_nl = MUX_s_1_2_2(or_1983_cse, mux_1394_nl, fsm_output[5]);
  assign mux_1400_nl = MUX_s_1_2_2(mux_1399_nl, mux_1395_nl, fsm_output[4]);
  assign and_dcpl_618 = ~(mux_1400_nl | (fsm_output[8]));
  assign and_dcpl_619 = and_dcpl_241 & and_dcpl_256;
  assign or_tmp_1203 = (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[2]) |
      (~ (fsm_output[4]));
  assign mux_1405_nl = MUX_s_1_2_2(or_tmp_1203, or_tmp_767, fsm_output[5]);
  assign or_2309_nl = (fsm_output[3]) | mux_1405_nl;
  assign or_1049_nl = (~ (fsm_output[2])) | (fsm_output[5]) | (fsm_output[4]);
  assign mux_1404_nl = MUX_s_1_2_2(or_1049_nl, or_349_cse, fsm_output[3]);
  assign mux_1406_nl = MUX_s_1_2_2(or_2309_nl, mux_1404_nl, fsm_output[6]);
  assign and_dcpl_620 = (~ mux_1406_nl) & and_dcpl_295;
  assign or_2322_nl = (fsm_output[5]) | or_tmp_728;
  assign mux_tmp_1421 = MUX_s_1_2_2(or_2699_cse, or_2322_nl, fsm_output[3]);
  assign or_tmp_1218 = (fsm_output[6]) | mux_tmp_1421;
  assign and_1303_nl = (fsm_output[2]) & (fsm_output[5]) & (fsm_output[4]);
  assign mux_1422_nl = MUX_s_1_2_2(and_1303_nl, and_1762_cse, fsm_output[3]);
  assign not_tmp_650 = ~((fsm_output[6]) | mux_1422_nl);
  assign mux_1424_nl = MUX_s_1_2_2(not_tmp_650, or_tmp_1132, fsm_output[7]);
  assign mux_1423_nl = MUX_s_1_2_2(not_tmp_650, or_tmp_1218, fsm_output[7]);
  assign mux_1425_nl = MUX_s_1_2_2(mux_1424_nl, mux_1423_nl, reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign and_dcpl_622 = ~(mux_1425_nl | (fsm_output[8]));
  assign and_dcpl_625 = (~((fsm_output[8]) | (fsm_output[0]) | (fsm_output[5])))
      & and_dcpl_45;
  assign or_tmp_1221 = (fsm_output[1]) | (fsm_output[2]) | (~ (fsm_output[4]));
  assign mux_tmp_1426 = MUX_s_1_2_2(or_tmp_1221, or_tmp_1128, fsm_output[3]);
  assign or_2328_nl = (fsm_output[4:1]!=4'b1000);
  assign mux_1427_nl = MUX_s_1_2_2(or_2328_nl, mux_tmp_1426, reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign and_dcpl_626 = (~ mux_1427_nl) & and_dcpl_625;
  assign and_dcpl_628 = and_dcpl_201 & (fsm_output[5]);
  assign mux_1435_nl = MUX_s_1_2_2((~ and_1559_cse), or_3185_cse, fsm_output[3]);
  assign nor_938_nl = ~((fsm_output[6]) | mux_1435_nl);
  assign nor_939_nl = ~((~ (fsm_output[6])) | (fsm_output[3]) | (~ and_1637_cse));
  assign mux_1436_nl = MUX_s_1_2_2(nor_938_nl, nor_939_nl, fsm_output[7]);
  assign and_dcpl_629 = mux_1436_nl & and_dcpl_628;
  assign mux_tmp_1440 = MUX_s_1_2_2((~ and_1637_cse), or_3185_cse, fsm_output[3]);
  assign mux_1449_nl = MUX_s_1_2_2(and_dcpl_383, and_1559_cse, fsm_output[0]);
  assign mux_1450_nl = MUX_s_1_2_2((~ or_3185_cse), mux_1449_nl, fsm_output[3]);
  assign and_dcpl_635 = mux_1450_nl & (~ (fsm_output[8])) & (~ (fsm_output[4])) &
      (fsm_output[5]) & and_dcpl_45;
  assign and_tmp_42 = (fsm_output[5]) & ((~((fsm_output[2:0]!=3'b101))) | (fsm_output[4]));
  assign mux_tmp_1451 = MUX_s_1_2_2(or_255_cse, or_270_cse, or_1732_cse);
  assign and_dcpl_641 = and_1474_cse & (fsm_output[5]);
  assign and_dcpl_642 = and_dcpl_641 & and_dcpl_420;
  assign or_dcpl_1108 = or_241_cse | or_dcpl_79;
  assign or_2395_cse = (fsm_output[5]) | (fsm_output[2]) | (fsm_output[4]);
  assign mux_tmp_1489 = MUX_s_1_2_2(or_2699_cse, or_2395_cse, fsm_output[3]);
  assign or_dcpl_1109 = (~ (fsm_output[5])) | (fsm_output[3]);
  assign or_dcpl_1114 = or_241_cse | or_dcpl_68;
  assign and_dcpl_650 = (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2])) & (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]);
  assign and_dcpl_651 = and_dcpl_650 & (~ reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1);
  assign or_dcpl_1116 = or_241_cse | or_dcpl_60;
  assign and_dcpl_656 = and_dcpl_650 & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1;
  assign or_dcpl_1118 = or_241_cse | or_dcpl_45;
  assign or_dcpl_1119 = (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b01);
  assign or_dcpl_1120 = or_dcpl_1119 | or_dcpl_79;
  assign or_dcpl_1121 = or_dcpl_1119 | or_dcpl_68;
  assign or_dcpl_1122 = or_dcpl_1119 | or_dcpl_60;
  assign or_dcpl_1123 = or_dcpl_1119 | or_dcpl_45;
  assign or_dcpl_1125 = or_dcpl_672 | or_dcpl_79;
  assign or_dcpl_1126 = or_dcpl_672 | or_dcpl_68;
  assign or_dcpl_1127 = or_dcpl_672 | or_dcpl_60;
  assign or_dcpl_1128 = or_dcpl_672 | or_dcpl_45;
  assign or_dcpl_1130 = or_dcpl_47 | or_dcpl_79;
  assign or_dcpl_1131 = or_dcpl_47 | or_dcpl_68;
  assign or_dcpl_1132 = or_dcpl_47 | or_dcpl_60;
  assign or_dcpl_1133 = or_dcpl_47 | or_dcpl_45;
  assign or_tmp_1291 = (fsm_output[7:4]!=4'b1000);
  assign or_tmp_1296 = (fsm_output[2]) | (~ (fsm_output[3])) | (fsm_output[4]) |
      (~ (fsm_output[7])) | (fsm_output[6]) | (fsm_output[8]);
  assign and_dcpl_718 = and_dcpl_307 & (fsm_output[7]);
  assign or_tmp_1316 = (~((fsm_output[4:3]!=2'b01))) | (fsm_output[8:6]!=3'b010);
  assign mux_tmp_1519 = MUX_s_1_2_2(or_tmp_507, or_tmp_812, fsm_output[4]);
  assign or_tmp_1320 = (fsm_output[3]) | (fsm_output[4]) | (~ (fsm_output[7])) |
      (~ (fsm_output[6])) | (fsm_output[8]);
  assign and_dcpl_721 = and_dcpl_591 & and_dcpl_335;
  assign mux_137_nl = MUX_s_1_2_2(or_2699_cse, or_349_cse, fsm_output[3]);
  assign not_tmp_699 = ~((fsm_output[6]) & mux_137_nl);
  assign and_dcpl_725 = and_dcpl_315 & and_dcpl_256;
  assign and_dcpl_726 = and_dcpl_376 & and_dcpl_256;
  assign or_dcpl_1134 = (fsm_output[5]) | (~ (fsm_output[3]));
  assign or_dcpl_1137 = nand_143_cse | or_dcpl_1077;
  assign or_dcpl_1138 = or_dcpl_1070 | or_750_cse;
  assign or_dcpl_1140 = (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1)
      | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd;
  assign or_dcpl_1141 = or_dcpl_1140 | or_dcpl_351;
  assign and_dcpl_727 = (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd)
      & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[1]);
  assign and_dcpl_728 = and_dcpl_727 & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]);
  assign and_dcpl_729 = and_dcpl_57 & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  assign and_dcpl_730 = and_dcpl_729 & and_dcpl_728;
  assign and_dcpl_731 = and_dcpl_61 & and_dcpl_383;
  assign and_dcpl_732 = and_dcpl_731 & and_dcpl_553;
  assign mux_tmp_1548 = MUX_s_1_2_2(mux_tmp_121, or_tmp_464, fsm_output[5]);
  assign mux_tmp_1549 = MUX_s_1_2_2(or_tmp_464, mux_tmp_121, fsm_output[5]);
  assign nand_tmp_66 = ~((fsm_output[5]) & (~ mux_tmp_121));
  assign and_dcpl_735 = and_dcpl_61 & and_1559_cse;
  assign and_dcpl_736 = and_dcpl_735 & and_dcpl_357 & (fsm_output[3]);
  assign and_dcpl_739 = and_dcpl_263 & nor_777_cse & and_dcpl_261;
  assign and_dcpl_740 = nor_973_cse & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  assign and_dcpl_743 = nor_tmp_99 & and_dcpl_383 & and_dcpl_553;
  assign and_dcpl_745 = nor_1026_cse & (fsm_output[3]);
  assign and_dcpl_747 = (~ (fsm_output[4])) & (fsm_output[2]) & (fsm_output[1]);
  assign and_dcpl_748 = and_dcpl_747 & and_dcpl_745;
  assign mux_tmp_1562 = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), fsm_output[7]);
  assign and_dcpl_751 = and_dcpl_45 & (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[1]);
  assign and_dcpl_753 = and_dcpl_735 & and_dcpl_745;
  assign and_dcpl_754 = and_dcpl_753 & and_dcpl_751 & and_dcpl_656;
  assign and_dcpl_758 = and_dcpl_45 & (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[1]));
  assign and_dcpl_760 = and_dcpl_753 & and_dcpl_758 & and_dcpl_512;
  assign and_dcpl_764 = and_dcpl_753 & and_dcpl_751 & and_dcpl_651;
  assign and_dcpl_768 = and_dcpl_753 & and_dcpl_758 & and_dcpl_525;
  assign and_dcpl_772 = and_dcpl_753 & and_dcpl_751 & and_dcpl_458;
  assign and_dcpl_776 = and_dcpl_753 & and_dcpl_758 & and_dcpl_468;
  assign and_dcpl_780 = and_dcpl_753 & and_dcpl_751 & and_dcpl_354;
  assign and_dcpl_784 = and_dcpl_753 & and_dcpl_758 & and_dcpl_539;
  assign and_dcpl_788 = and_dcpl_753 & and_dcpl_751 & and_dcpl_512;
  assign and_dcpl_792 = and_dcpl_753 & and_dcpl_751 & and_dcpl_525;
  assign and_dcpl_796 = and_dcpl_753 & and_dcpl_758 & and_dcpl_458;
  assign and_dcpl_800 = and_dcpl_753 & and_dcpl_751 & and_dcpl_468;
  assign and_dcpl_804 = and_dcpl_753 & and_dcpl_758 & and_dcpl_354;
  assign and_dcpl_810 = and_dcpl_181 & (~ (fsm_output[6]));
  assign and_dcpl_812 = and_dcpl_376 & and_dcpl_810 & (fsm_output[7]) & (LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1[4]);
  assign and_dcpl_813 = and_dcpl_231 & (~ (fsm_output[7]));
  assign and_dcpl_814 = and_dcpl_747 & and_dcpl_813;
  assign mux_tmp_1578 = MUX_s_1_2_2((~ (fsm_output[0])), (fsm_output[0]), fsm_output[5]);
  assign and_dcpl_817 = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & (~
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[1]));
  assign and_dcpl_818 = and_dcpl_817 & (~ (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]));
  assign and_dcpl_819 = and_dcpl_57 & (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1);
  assign and_dcpl_820 = and_dcpl_819 & and_dcpl_818;
  assign and_dcpl_821 = and_dcpl_736 & and_dcpl_820;
  assign or_tmp_1354 = (fsm_output[5]) | (fsm_output[0]);
  assign and_dcpl_825 = and_dcpl_727 & (~ (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]));
  assign and_dcpl_826 = and_dcpl_729 & and_dcpl_825;
  assign and_dcpl_827 = and_dcpl_736 & and_dcpl_826;
  assign and_dcpl_830 = and_dcpl_817 & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]);
  assign and_dcpl_831 = and_dcpl_819 & and_dcpl_830;
  assign and_dcpl_832 = and_dcpl_736 & and_dcpl_831;
  assign and_dcpl_835 = and_dcpl_549 & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]);
  assign and_dcpl_836 = and_dcpl_729 & and_dcpl_835;
  assign and_dcpl_837 = and_dcpl_736 & and_dcpl_836;
  assign and_dcpl_840 = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[1]);
  assign and_dcpl_841 = and_dcpl_840 & (~ (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]));
  assign and_dcpl_842 = and_dcpl_819 & and_dcpl_841;
  assign and_dcpl_843 = and_dcpl_736 & and_dcpl_842;
  assign or_2500_cse = (fsm_output[1]) | RESHAPE_2D_TO_3D_LOOP_2_2_and_cse;
  assign and_dcpl_847 = and_dcpl_205 & or_2500_cse & nor_1026_cse & (~ (fsm_output[3]))
      & and_dcpl_45;
  assign and_dcpl_850 = and_dcpl_729 & and_dcpl_550;
  assign and_dcpl_851 = and_dcpl_736 & and_dcpl_850;
  assign and_dcpl_854 = and_dcpl_840 & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]);
  assign and_dcpl_855 = and_dcpl_819 & and_dcpl_854;
  assign and_dcpl_856 = and_dcpl_736 & and_dcpl_855;
  assign and_dcpl_859 = and_dcpl_729 & and_dcpl_818;
  assign and_dcpl_860 = and_dcpl_736 & and_dcpl_859;
  assign and_dcpl_863 = and_dcpl_729 & and_dcpl_830;
  assign and_dcpl_864 = and_dcpl_736 & and_dcpl_863;
  assign and_dcpl_867 = and_dcpl_819 & and_dcpl_835;
  assign and_dcpl_868 = and_dcpl_736 & and_dcpl_867;
  assign and_dcpl_871 = and_dcpl_729 & and_dcpl_841;
  assign and_dcpl_872 = and_dcpl_736 & and_dcpl_871;
  assign and_dcpl_875 = and_dcpl_819 & and_dcpl_550;
  assign and_dcpl_876 = and_dcpl_736 & and_dcpl_875;
  assign and_dcpl_879 = and_dcpl_729 & and_dcpl_854;
  assign and_dcpl_880 = and_dcpl_736 & and_dcpl_879;
  assign and_dcpl_885 = (~ (fsm_output[5])) & (fsm_output[7]);
  assign or_tmp_1392 = ~((fsm_output[3]) & (fsm_output[0]) & (fsm_output[1]) & (~
      (fsm_output[4])));
  assign and_dcpl_888 = and_dcpl_731 & and_dcpl_256;
  assign and_dcpl_959 = and_dcpl_753 & and_dcpl_758 & and_dcpl_656;
  assign nor_946_nl = ~((or_2792_cse & (fsm_output[2])) | (fsm_output[4]));
  assign mux_1942_nl = MUX_s_1_2_2(nor_946_nl, or_tmp_728, fsm_output[5]);
  assign mux_tmp_1943 = MUX_s_1_2_2(mux_tmp_91, mux_1942_nl, fsm_output[3]);
  assign mux_1944_nl = MUX_s_1_2_2(nor_992_cse, or_tmp_728, fsm_output[5]);
  assign mux_tmp_1945 = MUX_s_1_2_2(mux_tmp_91, mux_1944_nl, fsm_output[3]);
  assign and_dcpl_983 = and_dcpl_376 & and_dcpl_810 & (fsm_output[7]) & (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign and_dcpl_987 = and_dcpl_819 & and_dcpl_825;
  assign and_dcpl_989 = and_dcpl_736 & and_dcpl_987;
  assign and_dcpl_999 = and_dcpl_753 & and_dcpl_758 & and_dcpl_651;
  assign and_dcpl_1000 = and_dcpl_819 & and_dcpl_728;
  assign mux_tmp_1990 = MUX_s_1_2_2(mux_806_cse, or_1983_cse, fsm_output[5]);
  assign mux_tmp_1993 = MUX_s_1_2_2(or_2249_cse, or_1983_cse, fsm_output[5]);
  assign and_dcpl_1003 = and_dcpl_736 & and_dcpl_1000;
  assign or_dcpl_1145 = or_76_cse | or_dcpl_1003;
  assign mux_tmp_2013 = MUX_s_1_2_2(or_1985_cse, or_tmp_914, fsm_output[4]);
  assign mux_tmp_2015 = MUX_s_1_2_2(or_1985_cse, or_2717_cse, fsm_output[4]);
  assign or_dcpl_1146 = or_dcpl_1022 | or_dcpl_1029;
  assign or_2744_nl = RESHAPE_2D_TO_3D_LOOP_2_2_and_cse | (fsm_output[1]) | (fsm_output[2])
      | (~ (fsm_output[4]));
  assign mux_tmp_2034 = MUX_s_1_2_2(or_2744_nl, or_tmp_1128, fsm_output[3]);
  assign or_2746_nl = (fsm_output[3]) | RESHAPE_2D_TO_3D_LOOP_2_2_and_cse | (fsm_output[1])
      | (fsm_output[2]) | (~ (fsm_output[4]));
  assign mux_2035_nl = MUX_s_1_2_2(or_2746_nl, mux_tmp_2034, reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign and_dcpl_1011 = (~ mux_2035_nl) & and_dcpl_625;
  assign and_dcpl_1033 = and_dcpl_376 & and_dcpl_810 & (fsm_output[7]) & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign and_dcpl_1034 = and_dcpl_362 & and_dcpl_199;
  assign mux_2066_nl = MUX_s_1_2_2((~ (fsm_output[4])), mux_tmp_1113, fsm_output[0]);
  assign mux_tmp_2067 = MUX_s_1_2_2(mux_2066_nl, or_tmp_330, fsm_output[3]);
  assign and_dcpl_1055 = (~(and_1559_cse & (fsm_output[0]))) & and_dcpl_201 & and_dcpl_199;
  assign and_dcpl_1061 = and_dcpl_735 & and_dcpl_553;
  assign or_tmp_1632 = and_1474_cse | (fsm_output[2]) | (fsm_output[4]);
  assign or_2784_nl = (fsm_output[5]) | or_tmp_1632;
  assign mux_2085_nl = MUX_s_1_2_2(or_2699_cse, or_2784_nl, fsm_output[3]);
  assign not_tmp_874 = ~((fsm_output[6]) & mux_2085_nl);
  assign or_tmp_1643 = (~ (fsm_output[4])) | (fsm_output[7]) | (fsm_output[6]) |
      (~ (fsm_output[8]));
  assign or_dcpl_1152 = nand_129_cse | or_dcpl_351;
  assign or_dcpl_1155 = or_dcpl_377 | or_dcpl_332;
  assign or_dcpl_1156 = nand_129_cse | or_dcpl_337;
  assign or_dcpl_1158 = or_dcpl_377 | or_dcpl_342;
  assign or_dcpl_1159 = nand_129_cse | or_dcpl_342;
  assign or_dcpl_1160 = or_dcpl_377 | or_dcpl_337;
  assign or_dcpl_1161 = nand_129_cse | or_dcpl_332;
  assign or_dcpl_1162 = or_dcpl_377 | or_dcpl_351;
  assign or_dcpl_1163 = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 |
      (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd);
  assign or_dcpl_1164 = or_dcpl_1163 | or_dcpl_351;
  assign or_dcpl_1165 = or_dcpl_1140 | or_dcpl_332;
  assign or_dcpl_1166 = or_dcpl_1163 | or_dcpl_337;
  assign or_dcpl_1167 = or_dcpl_1140 | or_dcpl_342;
  assign or_dcpl_1168 = or_dcpl_1163 | or_dcpl_342;
  assign or_dcpl_1169 = or_dcpl_1140 | or_dcpl_337;
  assign or_dcpl_1170 = or_dcpl_1163 | or_dcpl_332;
  assign and_dcpl_1073 = (~ mux_tmp_2034) & and_dcpl_625;
  assign and_dcpl_1082 = and_dcpl_211 & (fsm_output[5]) & and_dcpl_813;
  assign and_dcpl_1084 = or_dcpl_1138 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1088 = or_dcpl_1084 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1091 = or_dcpl_1071 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1094 = or_dcpl_1092 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1097 = or_dcpl_1090 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1100 = or_dcpl_1088 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1103 = or_dcpl_1086 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1106 = or_dcpl_1079 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1109 = or_dcpl_1067 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1112 = or_dcpl_1087 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1115 = or_dcpl_1089 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1118 = or_dcpl_1091 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1121 = or_dcpl_1073 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1124 = or_dcpl_1083 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1127 = or_dcpl_1085 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1130 = or_dcpl_1137 & and_dcpl_191 & and_dcpl_1082;
  assign and_dcpl_1141 = and_dcpl_243 & (fsm_output[7]);
  assign and_dcpl_1145 = and_dcpl_279 & and_dcpl_45;
  assign or_2834_cse = (fsm_output[6:5]!=2'b01);
  assign nor_953_nl = ~(nor_777_cse | (fsm_output[6:5]!=2'b01));
  assign nor_954_nl = ~((fsm_output[1]) | (fsm_output[0]) | (fsm_output[5]) | (~
      (fsm_output[6])));
  assign mux_2111_nl = MUX_s_1_2_2(nor_953_nl, nor_954_nl, fsm_output[3]);
  assign or_2833_nl = (fsm_output[6:5]!=2'b10);
  assign mux_2110_nl = MUX_s_1_2_2(or_2834_cse, or_2833_nl, or_1732_cse);
  assign nor_955_nl = ~((fsm_output[3]) | mux_2110_nl);
  assign mux_2112_nl = MUX_s_1_2_2(mux_2111_nl, nor_955_nl, fsm_output[2]);
  assign nor_956_nl = ~((fsm_output[2]) | (fsm_output[3]) | (fsm_output[1]) | (~
      (fsm_output[0])) | (fsm_output[5]) | (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1)
      | (fsm_output[6]));
  assign mux_2113_nl = MUX_s_1_2_2(mux_2112_nl, nor_956_nl, fsm_output[4]);
  assign and_dcpl_1151 = mux_2113_nl & and_dcpl_295;
  assign and_dcpl_1152 = and_dcpl_186 & and_dcpl_190;
  assign or_tmp_1664 = (fsm_output[8:5]!=4'b1001);
  assign mux_2115_nl = MUX_s_1_2_2(or_tmp_507, or_1197_cse, fsm_output[5]);
  assign mux_tmp_2116 = MUX_s_1_2_2(mux_2115_nl, or_tmp_1664, fsm_output[4]);
  assign nor_957_nl = ~((~ (fsm_output[8])) | (fsm_output[6]));
  assign mux_2117_nl = MUX_s_1_2_2(nor_957_nl, and_dcpl_307, fsm_output[7]);
  assign nand_tmp_99 = ~((fsm_output[5]) & mux_2117_nl);
  assign mux_2118_nl = MUX_s_1_2_2(nand_tmp_99, or_tmp_1664, fsm_output[4]);
  assign mux_tmp_2119 = MUX_s_1_2_2(mux_2118_nl, mux_tmp_2116, fsm_output[2]);
  assign or_tmp_1671 = nor_646_cse | (fsm_output[8:6]!=3'b100);
  assign mux_tmp_2121 = MUX_s_1_2_2(mux_tmp_2119, or_tmp_1671, fsm_output[3]);
  assign and_dcpl_1154 = and_dcpl_449 & and_1474_cse & and_dcpl_261;
  assign and_dcpl_1162 = and_dcpl_241 & and_dcpl_198 & (~ (z_out_5[2])) & and_dcpl_148;
  assign or_tmp_1690 = (~ (fsm_output[1])) | (~ (fsm_output[7])) | (fsm_output[8]);
  assign mux_2149_nl = MUX_s_1_2_2(or_822_cse, mux_623_cse, nor_354_cse);
  assign mux_2147_nl = MUX_s_1_2_2(mux_623_cse, or_822_cse, and_1474_cse);
  assign nand_286_nl = ~((fsm_output[0]) & (fsm_output[1]) & (fsm_output[7]) & (~
      (fsm_output[8])));
  assign mux_2148_nl = MUX_s_1_2_2(mux_2147_nl, nand_286_nl, fsm_output[3]);
  assign mux_2150_nl = MUX_s_1_2_2(mux_2149_nl, mux_2148_nl, fsm_output[2]);
  assign mux_2151_nl = MUX_s_1_2_2(or_822_cse, mux_2150_nl, fsm_output[4]);
  assign nand_101_nl = ~((fsm_output[3]) & (~(nor_777_cse | (fsm_output[8:7]!=2'b01))));
  assign or_2868_nl = (fsm_output[1]) | (~ (fsm_output[7])) | (fsm_output[8]);
  assign mux_2144_nl = MUX_s_1_2_2(or_tmp_1690, or_2868_nl, fsm_output[0]);
  assign or_2869_nl = (fsm_output[3]) | mux_2144_nl;
  assign mux_2145_nl = MUX_s_1_2_2(nand_101_nl, or_2869_nl, fsm_output[2]);
  assign or_2872_nl = (fsm_output[4]) | mux_2145_nl;
  assign mux_2152_nl = MUX_s_1_2_2(mux_2151_nl, or_2872_nl, fsm_output[5]);
  assign or_2866_nl = nor_355_cse | (fsm_output[8:7]!=2'b01);
  assign mux_2142_nl = MUX_s_1_2_2(or_tmp_1690, or_2866_nl, fsm_output[3]);
  assign mux_2143_nl = MUX_s_1_2_2(mux_2142_nl, or_361_cse, or_2395_cse);
  assign mux_tmp_2153 = MUX_s_1_2_2(mux_2152_nl, mux_2143_nl, fsm_output[6]);
  assign or_dcpl_1178 = or_dcpl_770 | nand_163_cse;
  assign nor_964_cse = ~((fsm_output[1]) | (fsm_output[4]));
  assign mux_2172_nl = MUX_s_1_2_2(or_1197_cse, mux_tmp_604, fsm_output[4]);
  assign mux_2171_nl = MUX_s_1_2_2(mux_tmp_604, mux_624_cse, fsm_output[4]);
  assign mux_2173_nl = MUX_s_1_2_2(mux_2172_nl, mux_2171_nl, fsm_output[1]);
  assign or_2901_nl = (fsm_output[1:0]!=2'b10) | (~ (z_out_5[2])) | (fsm_output[4]);
  assign mux_2170_nl = MUX_s_1_2_2(or_1197_cse, mux_tmp_604, or_2901_nl);
  assign mux_2174_nl = MUX_s_1_2_2(mux_2173_nl, mux_2170_nl, fsm_output[3]);
  assign and_1544_nl = nand_197_cse & (fsm_output[4]);
  assign mux_2168_nl = MUX_s_1_2_2(mux_tmp_604, mux_624_cse, and_1544_nl);
  assign mux_2164_nl = MUX_s_1_2_2(mux_tmp_604, or_tmp_507, fsm_output[4]);
  assign mux_2162_nl = MUX_s_1_2_2(or_822_cse, or_361_cse, or_1879_cse);
  assign mux_2165_nl = MUX_s_1_2_2(mux_2164_nl, mux_2162_nl, and_1474_cse);
  assign mux_2169_nl = MUX_s_1_2_2(mux_2168_nl, mux_2165_nl, fsm_output[3]);
  assign mux_2175_nl = MUX_s_1_2_2(mux_2174_nl, mux_2169_nl, fsm_output[2]);
  assign or_2897_nl = (~((~((~ (fsm_output[1])) | (fsm_output[4]))) | (fsm_output[6])))
      | (fsm_output[8:7]!=2'b01);
  assign or_2894_nl = (~(nor_964_cse | (fsm_output[6]))) | (fsm_output[8:7]!=2'b01);
  assign mux_2160_nl = MUX_s_1_2_2(or_2897_nl, or_2894_nl, fsm_output[0]);
  assign or_2890_nl = (fsm_output[3:2]!=2'b01);
  assign mux_2161_nl = MUX_s_1_2_2(mux_2160_nl, or_tmp_507, or_2890_nl);
  assign mux_tmp_2176 = MUX_s_1_2_2(mux_2175_nl, mux_2161_nl, fsm_output[5]);
  assign or_dcpl_1180 = or_dcpl_794 | or_1435_cse;
  assign or_dcpl_1181 = or_dcpl_770 | or_1431_cse;
  assign or_dcpl_1183 = or_dcpl_770 | or_1420_cse;
  assign or_dcpl_1184 = or_dcpl_794 | or_1420_cse;
  assign or_dcpl_1186 = or_dcpl_791 | or_1435_cse;
  assign or_dcpl_1187 = or_dcpl_774 | nand_163_cse;
  assign or_dcpl_1188 = or_dcpl_774 | or_1435_cse;
  assign or_dcpl_1189 = or_dcpl_791 | or_1420_cse;
  assign and_dcpl_1193 = and_dcpl_376 & and_dcpl_190;
  assign and_dcpl_1194 = and_dcpl_239 & and_dcpl_190;
  assign and_dcpl_1195 = and_dcpl_186 & and_dcpl_293;
  assign or_dcpl_1195 = ~((z_out_11[0]) & (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[0]));
  assign or_dcpl_1196 = (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2:1]!=2'b10);
  assign or_dcpl_1198 = (z_out_11[0]) | (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[0]);
  assign or_dcpl_1199 = (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2:1]!=2'b00);
  assign or_dcpl_1201 = (z_out_11[0]) | (~ (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[0]));
  assign or_dcpl_1203 = (~ (z_out_11[0])) | (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[0]);
  assign or_dcpl_1209 = (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2:1]!=2'b01);
  assign and_dcpl_1199 = and_dcpl_241 & and_dcpl_221;
  assign and_1546_nl = (fsm_output[5]) & (fsm_output[2]) & (fsm_output[4]) & (~ (fsm_output[8]));
  assign nor_968_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_2251_nl = MUX_s_1_2_2(and_1546_nl, nor_968_nl, fsm_output[3]);
  assign nand_tmp_104 = ~((fsm_output[6]) & mux_2251_nl);
  assign or_3055_nl = (fsm_output[6]) | (~((~((fsm_output[5:0]==6'b111111))) & (fsm_output[8])));
  assign mux_tmp_2252 = MUX_s_1_2_2(or_3055_nl, nand_tmp_104, fsm_output[7]);
  assign or_1418_nl = (fsm_output[2:0]!=3'b011);
  assign mux_2253_nl = MUX_s_1_2_2(and_dcpl_252, (fsm_output[8]), or_1418_nl);
  assign nand_295_nl = ~(nand_240_cse & (fsm_output[8]));
  assign mux_2254_nl = MUX_s_1_2_2((~ mux_2253_nl), nand_295_nl, fsm_output[5]);
  assign mux_2255_nl = MUX_s_1_2_2((~ (fsm_output[8])), mux_2254_nl, fsm_output[3]);
  assign or_3058_nl = (fsm_output[6]) | mux_2255_nl;
  assign mux_2256_itm = MUX_s_1_2_2(or_3058_nl, nand_tmp_104, fsm_output[7]);
  assign and_dcpl_1225 = and_dcpl_263 & and_dcpl_211 & and_dcpl_275;
  assign and_dcpl_1227 = and_dcpl_263 & and_dcpl_200 & and_dcpl_261;
  assign and_1550_nl = (fsm_output[5:0]==6'b111111);
  assign nor_969_nl = ~((fsm_output[5:0]!=6'b000000));
  assign mux_2259_nl = MUX_s_1_2_2(and_1550_nl, nor_969_nl, fsm_output[6]);
  assign and_dcpl_1232 = mux_2259_nl & (fsm_output[8:7]==2'b10);
  assign mux_868_nl = MUX_s_1_2_2(or_dcpl_1050, nor_tmp_282, fsm_output[5]);
  assign mux_869_nl = MUX_s_1_2_2(mux_868_nl, mux_tmp_91, fsm_output[3]);
  assign rms_norm_16_div_cmp_a_mx0c0 = (~ mux_869_nl) & and_dcpl_308;
  assign attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c0 = and_dcpl_342 &
      and_dcpl_336 & and_dcpl_335;
  assign attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c9 = and_dcpl_360 &
      and_dcpl_355 & and_dcpl_354;
  assign nor_998_cse = ~(nor_777_cse | (fsm_output[4]));
  assign nor_999_nl = ~((~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[4])
      | (fsm_output[8]));
  assign mux_1007_nl = MUX_s_1_2_2(nor_999_nl, (fsm_output[8]), fsm_output[5]);
  assign mux_1008_nl = MUX_s_1_2_2((~ mux_1007_nl), mux_958_cse, fsm_output[6]);
  assign nand_322_nl = ~(or_1732_cse & (fsm_output[4]) & (fsm_output[8]));
  assign nor_1001_nl = ~(nor_176_cse | (fsm_output[8]));
  assign mux_1005_nl = MUX_s_1_2_2(nand_322_nl, nor_1001_nl, fsm_output[5]);
  assign or_1952_nl = nor_964_cse | (fsm_output[8]);
  assign or_1950_nl = (~((~ LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4) | (~ (fsm_output[1]))
      | (fsm_output[4]))) | (fsm_output[8]);
  assign mux_1003_nl = MUX_s_1_2_2(or_1952_nl, or_1950_nl, fsm_output[0]);
  assign mux_1004_nl = MUX_s_1_2_2(mux_1003_nl, or_133_cse, fsm_output[5]);
  assign mux_1006_nl = MUX_s_1_2_2(mux_1005_nl, mux_1004_nl, fsm_output[6]);
  assign mux_1009_nl = MUX_s_1_2_2(mux_1008_nl, mux_1006_nl, fsm_output[3]);
  assign nand_323_nl = ~((fsm_output[5]) & ((or_1732_cse & (fsm_output[4])) | (fsm_output[8])));
  assign mux_1001_nl = MUX_s_1_2_2(nand_323_nl, mux_958_cse, fsm_output[6]);
  assign nand_325_nl = ~(nand_263_cse & (fsm_output[8]));
  assign mux_998_nl = MUX_s_1_2_2(or_dcpl_959, nand_325_nl, fsm_output[5]);
  assign or_1944_nl = (fsm_output[1]) | (fsm_output[4]) | (fsm_output[8]);
  assign mux_997_nl = MUX_s_1_2_2((fsm_output[8]), or_1944_nl, fsm_output[5]);
  assign mux_999_nl = MUX_s_1_2_2(mux_998_nl, mux_997_nl, fsm_output[6]);
  assign mux_1002_nl = MUX_s_1_2_2(mux_1001_nl, mux_999_nl, fsm_output[3]);
  assign mux_1010_nl = MUX_s_1_2_2(mux_1009_nl, mux_1002_nl, fsm_output[2]);
  assign mux_993_nl = MUX_s_1_2_2(or_tmp_878, (fsm_output[8]), fsm_output[5]);
  assign or_1943_nl = (fsm_output[5]) | (fsm_output[1]) | (fsm_output[4]) | (fsm_output[8]);
  assign mux_994_nl = MUX_s_1_2_2(mux_993_nl, or_1943_nl, fsm_output[6]);
  assign mux_991_nl = MUX_s_1_2_2(or_tmp_878, or_tmp_48, fsm_output[5]);
  assign or_1940_nl = (~ (fsm_output[5])) | (fsm_output[0]) | (fsm_output[1]) | (~
      (fsm_output[4])) | (fsm_output[8]);
  assign mux_992_nl = MUX_s_1_2_2(mux_991_nl, or_1940_nl, fsm_output[6]);
  assign mux_995_nl = MUX_s_1_2_2(mux_994_nl, mux_992_nl, fsm_output[3]);
  assign or_1939_nl = (fsm_output[1]) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign or_1938_nl = (~ (fsm_output[1])) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_987_nl = MUX_s_1_2_2(or_1939_nl, or_1938_nl, fsm_output[0]);
  assign or_1937_nl = nor_998_cse | (fsm_output[8]);
  assign mux_988_nl = MUX_s_1_2_2(mux_987_nl, or_1937_nl, fsm_output[5]);
  assign or_1934_nl = (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_989_nl = MUX_s_1_2_2(mux_988_nl, or_1934_nl, fsm_output[6]);
  assign or_1932_nl = (fsm_output[0]) | (~ (fsm_output[1])) | (fsm_output[4]) | (fsm_output[8]);
  assign or_1931_nl = (~((fsm_output[0]) | (~ (fsm_output[1])) | (fsm_output[4])))
      | (fsm_output[8]);
  assign mux_986_nl = MUX_s_1_2_2(or_1932_nl, or_1931_nl, fsm_output[5]);
  assign or_1933_nl = (fsm_output[6]) | mux_986_nl;
  assign mux_990_nl = MUX_s_1_2_2(mux_989_nl, or_1933_nl, fsm_output[3]);
  assign mux_996_nl = MUX_s_1_2_2(mux_995_nl, mux_990_nl, fsm_output[2]);
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c0 = MUX_s_1_2_2(mux_1010_nl,
      mux_996_nl, fsm_output[7]);
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c2 = (~(((LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0==4'b1111)
      & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4) | mux_tmp_975)) & and_dcpl_202
      & (~ (fsm_output[1])) & (fsm_output[5]) & (~ (fsm_output[3]));
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c3 = (~(mux_tmp_975 | (fsm_output[8])))
      & and_1771_cse & (~ (fsm_output[1])) & and_dcpl_189 & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4
      & (LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0==4'b1111);
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c5 = and_dcpl_241 & and_dcpl_181
      & (fsm_output[6]) & (~((fsm_output[7]) | LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4));
  assign mux_1022_nl = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), fsm_output[5]);
  assign mux_1023_nl = MUX_s_1_2_2(mux_1022_nl, or_2834_cse, fsm_output[1]);
  assign nor_1019_nl = ~((fsm_output[3]) | mux_1023_nl);
  assign nor_1020_nl = ~((fsm_output[1]) | (~ (fsm_output[5])) | (fsm_output[6]));
  assign nor_1021_nl = ~((~ (fsm_output[3])) | (~ (fsm_output[5])) | (fsm_output[6]));
  assign mux_1021_nl = MUX_s_1_2_2(nor_1020_nl, nor_1021_nl, fsm_output[0]);
  assign mux_1024_nl = MUX_s_1_2_2(nor_1019_nl, mux_1021_nl, fsm_output[2]);
  assign nor_1022_nl = ~((~(and_1474_cse | (fsm_output[5]))) | (fsm_output[6]));
  assign nor_1023_nl = ~((~((~((fsm_output[3]) | (fsm_output[1]))) | (fsm_output[5])))
      | (fsm_output[6]));
  assign nor_1024_nl = ~((~(nor_354_cse | (fsm_output[5]))) | (fsm_output[6]));
  assign mux_1019_nl = MUX_s_1_2_2(nor_1023_nl, nor_1024_nl, fsm_output[0]);
  assign mux_1020_nl = MUX_s_1_2_2(nor_1022_nl, mux_1019_nl, fsm_output[2]);
  assign mux_1025_nl = MUX_s_1_2_2(mux_1024_nl, mux_1020_nl, fsm_output[4]);
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c7 = mux_1025_nl & and_dcpl_295;
  assign mux_1029_nl = MUX_s_1_2_2(or_tmp_728, or_tmp_704, fsm_output[0]);
  assign mux_1030_nl = MUX_s_1_2_2((~ mux_1029_nl), or_tmp_767, fsm_output[5]);
  assign mux_1031_nl = MUX_s_1_2_2(mux_tmp_91, mux_1030_nl, fsm_output[3]);
  assign nand_49_nl = ~((fsm_output[6]) & (~ mux_1031_nl));
  assign mux_1032_nl = MUX_s_1_2_2(nand_49_nl, or_tmp_913, fsm_output[7]);
  assign for_for_strm_in_tmp_sva_31_2_mx0c1 = ~(mux_1032_nl | (fsm_output[8]));
  assign GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c0 = and_dcpl_342 & and_dcpl_417 &
      and_dcpl_335;
  assign GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c1 = or_dcpl_1067 & and_dcpl_185 &
      and_dcpl_422;
  assign GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c2 = and_dcpl_289 & and_dcpl_425;
  assign GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c4 = and_dcpl_186 & and_dcpl_256;
  assign GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c7 = and_dcpl_192 & and_dcpl_293;
  assign GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c9 = and_dcpl_315 & and_dcpl_182;
  assign GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c10 = and_dcpl_327 & and_dcpl_291;
  assign attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c0 = and_dcpl_342 &
      and_dcpl_417 & and_dcpl_453;
  assign attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c1 = or_dcpl_1073 &
      and_dcpl_185 & and_dcpl_422;
  assign nor_1031_nl = ~((~((fsm_output[3:0]!=4'b0010))) | (fsm_output[8]));
  assign nand_330_nl = ~((~((fsm_output[3:2]==2'b11))) & (fsm_output[8]));
  assign mux_1078_nl = MUX_s_1_2_2(nor_1031_nl, nand_330_nl, fsm_output[4]);
  assign or_2029_cse = (fsm_output[6:5]!=2'b00) | mux_1078_nl;
  assign or_3163_cse = (z_out_5[2]) | (fsm_output[0]);
  assign nor_1032_nl = ~((fsm_output[3]) | (~ (fsm_output[0])) | (~ (fsm_output[1]))
      | (fsm_output[8]));
  assign nor_1033_nl = ~((fsm_output[3]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[8]));
  assign mux_1076_nl = MUX_s_1_2_2(nor_1032_nl, nor_1033_nl, fsm_output[2]);
  assign nand_50_cse = ~((~((fsm_output[5:4]!=2'b01))) & mux_1076_nl);
  assign or_2022_nl = (or_3163_cse & (fsm_output[1])) | (fsm_output[8]);
  assign mux_1073_nl = MUX_s_1_2_2(or_1848_cse, or_2022_nl, fsm_output[3]);
  assign mux_1074_cse = MUX_s_1_2_2(mux_1073_nl, (fsm_output[8]), or_255_cse);
  assign or_2019_nl = (~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b00) |
      (~ reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0])
      | (fsm_output[4:0]!=5'b10111))) | (fsm_output[8]);
  assign mux_1075_nl = MUX_s_1_2_2(mux_1074_cse, or_2019_nl, fsm_output[5]);
  assign mux_1077_nl = MUX_s_1_2_2(nand_50_cse, mux_1075_nl, fsm_output[6]);
  assign mux_1079_itm = MUX_s_1_2_2(or_2029_cse, mux_1077_nl, fsm_output[7]);
  assign mux_1088_nl = MUX_s_1_2_2(or_tmp_104, or_262_cse, fsm_output[0]);
  assign mux_1089_cse = MUX_s_1_2_2(mux_1088_nl, (fsm_output[8]), or_2797_cse);
  assign or_2038_nl = nor_355_cse | (fsm_output[8]);
  assign mux_1085_nl = MUX_s_1_2_2(or_262_cse, or_2038_nl, fsm_output[3]);
  assign mux_1086_nl = MUX_s_1_2_2(mux_1085_nl, (fsm_output[8]), fsm_output[4]);
  assign nand_52_nl = ~((fsm_output[7]) & (~ mux_1086_nl));
  assign mux_1087_cse = MUX_s_1_2_2(nand_52_nl, or_361_cse, fsm_output[5]);
  assign nand_332_nl = ~(nand_381_cse & (fsm_output[8]));
  assign nor_1035_nl = ~(and_1474_cse | (fsm_output[8]));
  assign nor_1036_nl = ~((~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[8]));
  assign mux_1081_nl = MUX_s_1_2_2(nor_1035_nl, nor_1036_nl, fsm_output[3]);
  assign nand_51_nl = ~((fsm_output[4]) & mux_1081_nl);
  assign mux_1082_nl = MUX_s_1_2_2(nand_332_nl, nand_51_nl, fsm_output[7]);
  assign mux_1080_nl = MUX_s_1_2_2(or_262_cse, or_tmp_104, fsm_output[0]);
  assign or_2034_nl = (~ (fsm_output[7])) | (fsm_output[4]) | (fsm_output[3]) | mux_1080_nl;
  assign mux_1083_nl = MUX_s_1_2_2(mux_1082_nl, or_2034_nl, fsm_output[5]);
  assign mux_1084_cse = MUX_s_1_2_2(mux_1083_nl, or_361_cse, fsm_output[6]);
  assign or_2039_nl = (~ (fsm_output[4])) | (fsm_output[3]) | (~ (fsm_output[0]))
      | (~ (fsm_output[1])) | (fsm_output[8]);
  assign mux_1090_nl = MUX_s_1_2_2((~ mux_1089_cse), or_2039_nl, fsm_output[7]);
  assign or_2041_nl = (fsm_output[5]) | mux_1090_nl;
  assign mux_1091_nl = MUX_s_1_2_2(or_2041_nl, mux_1087_cse, fsm_output[6]);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c7 = MUX_s_1_2_2(mux_1091_nl,
      mux_1084_cse, fsm_output[2]);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c9 = and_dcpl_360 &
      and_dcpl_355 & and_dcpl_458;
  assign attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c0 = and_dcpl_342 &
      and_dcpl_336 & and_dcpl_462;
  assign attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c1 = or_dcpl_1079 &
      and_dcpl_185 & and_dcpl_422;
  assign or_2068_nl = (~ (fsm_output[4])) | (fsm_output[3]) | (~ (fsm_output[1]))
      | (fsm_output[8]);
  assign mux_1110_nl = MUX_s_1_2_2((~ mux_1089_cse), or_2068_nl, fsm_output[7]);
  assign or_2070_nl = (fsm_output[5]) | mux_1110_nl;
  assign mux_1111_nl = MUX_s_1_2_2(or_2070_nl, mux_1087_cse, fsm_output[6]);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c7 = MUX_s_1_2_2(mux_1111_nl,
      mux_1084_cse, fsm_output[2]);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c9 = and_dcpl_360 &
      and_dcpl_355 & and_dcpl_468;
  assign apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c0 = and_dcpl_342 &
      and_dcpl_417 & and_dcpl_471;
  assign apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c1 = or_dcpl_1083 &
      and_dcpl_185 & and_dcpl_422;
  assign attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c0 = and_dcpl_342 & and_dcpl_417
      & and_dcpl_433;
  assign attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c1 = or_dcpl_1089 & and_dcpl_185
      & and_dcpl_422;
  assign mux_1129_nl = MUX_s_1_2_2(mux_1125_cse, mux_tmp_1120, fsm_output[0]);
  assign mux_1130_nl = MUX_s_1_2_2(mux_1122_cse, mux_1129_nl, fsm_output[2]);
  assign mux_1126_nl = MUX_s_1_2_2(or_1984_cse, mux_tmp_1120, fsm_output[4]);
  assign mux_1127_nl = MUX_s_1_2_2(mux_1126_nl, mux_1125_cse, fsm_output[0]);
  assign mux_1128_nl = MUX_s_1_2_2(mux_1127_nl, mux_tmp_1120, fsm_output[2]);
  assign mux_1131_nl = MUX_s_1_2_2(mux_1130_nl, mux_1128_nl, fsm_output[1]);
  assign mux_1121_nl = MUX_s_1_2_2(mux_tmp_1120, or_tmp_507, fsm_output[4]);
  assign mux_1123_nl = MUX_s_1_2_2(mux_1122_cse, mux_1121_nl, fsm_output[2]);
  assign mux_1132_cse = MUX_s_1_2_2(mux_1131_nl, mux_1123_nl, fsm_output[3]);
  assign attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c5 = and_dcpl_185 & ((fsm_output[1])
      ^ (fsm_output[3])) & and_dcpl_338 & and_dcpl_148;
  assign attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c8 = and_dcpl_350 & and_dcpl_182;
  assign attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c10 = and_dcpl_360 &
      and_dcpl_513 & and_dcpl_512;
  assign attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c0 = and_dcpl_342 & and_dcpl_336
      & and_dcpl_453;
  assign attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c1 = or_dcpl_1090 & and_dcpl_185
      & and_dcpl_422;
  assign or_2095_nl = ((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]==2'b11) & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1
      & (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0])) & (fsm_output[4:0]==5'b10111))
      | (fsm_output[8:6]!=3'b011);
  assign mux_1147_itm = MUX_s_1_2_2(mux_1132_cse, or_2095_nl, fsm_output[5]);
  assign attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c10 = and_dcpl_360 &
      and_dcpl_513 & and_dcpl_525;
  assign attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c0 = and_dcpl_342 & and_dcpl_417
      & and_dcpl_528;
  assign attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c1 = or_dcpl_1091 & and_dcpl_185
      & and_dcpl_422;
  assign or_2110_nl = ((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]==2'b11) & (~
      reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) & (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0])
      & (fsm_output[4:0]==5'b10111)) | (fsm_output[8:6]!=3'b011);
  assign mux_1177_itm = MUX_s_1_2_2(mux_1132_cse, or_2110_nl, fsm_output[5]);
  assign attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c10 = and_dcpl_360 &
      and_dcpl_513 & and_dcpl_468;
  assign attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c0 = and_dcpl_342 & and_dcpl_336
      & and_dcpl_528;
  assign attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c1 = or_dcpl_1092 & and_dcpl_185
      & and_dcpl_422;
  assign mux_1193_nl = MUX_s_1_2_2(or_1197_cse, mux_tmp_1183, fsm_output[4]);
  assign mux_1191_nl = MUX_s_1_2_2(or_1984_cse, mux_tmp_1187, fsm_output[4]);
  assign mux_1192_nl = MUX_s_1_2_2(mux_1191_nl, mux_tmp_1183, fsm_output[0]);
  assign mux_1194_nl = MUX_s_1_2_2(mux_1193_nl, mux_1192_nl, fsm_output[2]);
  assign mux_1188_nl = MUX_s_1_2_2(or_1197_cse, mux_tmp_1187, fsm_output[4]);
  assign mux_1189_nl = MUX_s_1_2_2(mux_tmp_1185, mux_1188_nl, fsm_output[0]);
  assign mux_1190_nl = MUX_s_1_2_2(mux_1189_nl, mux_tmp_1183, fsm_output[2]);
  assign mux_1195_nl = MUX_s_1_2_2(mux_1194_nl, mux_1190_nl, fsm_output[1]);
  assign mux_1184_nl = MUX_s_1_2_2(mux_tmp_1183, mux_tmp_1178, fsm_output[4]);
  assign mux_1186_nl = MUX_s_1_2_2(mux_tmp_1185, mux_1184_nl, fsm_output[2]);
  assign mux_1196_nl = MUX_s_1_2_2(mux_1195_nl, mux_1186_nl, fsm_output[3]);
  assign or_2121_nl = (fsm_output[4]) | mux_tmp_1178;
  assign and_1593_nl = (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]==2'b11) & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1
      & (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]);
  assign mux_1180_nl = MUX_s_1_2_2(mux_tmp_1179, or_2121_nl, and_1593_nl);
  assign mux_1181_nl = MUX_s_1_2_2(mux_tmp_1178, mux_1180_nl, and_1572_cse);
  assign mux_1182_nl = MUX_s_1_2_2(mux_1181_nl, mux_tmp_1179, fsm_output[3]);
  assign mux_1197_itm = MUX_s_1_2_2(mux_1196_nl, mux_1182_nl, fsm_output[5]);
  assign nor_1043_nl = ~((fsm_output[2]) | (fsm_output[1]) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[8]));
  assign and_1595_nl = (fsm_output[2]) & (fsm_output[3]) & (fsm_output[8]);
  assign mux_1205_nl = MUX_s_1_2_2(nor_1043_nl, and_1595_nl, fsm_output[4]);
  assign or_2130_nl = (or_2792_cse & (fsm_output[3])) | (fsm_output[8]);
  assign mux_1203_nl = MUX_s_1_2_2(or_2130_nl, or_tmp_1035, fsm_output[2]);
  assign mux_1204_nl = MUX_s_1_2_2((fsm_output[8]), mux_1203_nl, fsm_output[4]);
  assign mux_1206_nl = MUX_s_1_2_2(mux_1205_nl, mux_1204_nl, fsm_output[5]);
  assign or_2132_nl = (fsm_output[6]) | mux_1206_nl;
  assign or_2129_nl = (~ (fsm_output[1])) | (fsm_output[3]) | (fsm_output[8]);
  assign mux_1201_nl = MUX_s_1_2_2(or_2129_nl, or_tmp_1035, fsm_output[2]);
  assign or_3166_nl = (fsm_output[5:4]!=2'b01) | mux_1201_nl;
  assign or_2127_nl = (~ (fsm_output[3])) | (fsm_output[8]);
  assign or_2126_nl = (z_out_5[2]) | (~ (fsm_output[3])) | (fsm_output[8]);
  assign mux_1198_nl = MUX_s_1_2_2(or_2126_nl, (fsm_output[8]), fsm_output[0]);
  assign mux_1199_nl = MUX_s_1_2_2(or_2127_nl, mux_1198_nl, fsm_output[1]);
  assign mux_1200_nl = MUX_s_1_2_2(mux_1199_nl, (fsm_output[8]), or_2395_cse);
  assign mux_1202_nl = MUX_s_1_2_2(or_3166_nl, mux_1200_nl, fsm_output[6]);
  assign attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c10 = MUX_s_1_2_2(or_2132_nl,
      mux_1202_nl, fsm_output[7]);
  assign attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c12 = and_dcpl_360 &
      and_dcpl_513 & and_dcpl_539;
  assign or_2184_nl = and_1771_cse | (fsm_output[8]);
  assign mux_1270_nl = MUX_s_1_2_2(mux_tmp_967, or_2184_nl, fsm_output[1]);
  assign mux_1271_nl = MUX_s_1_2_2(mux_tmp_968, mux_1270_nl, fsm_output[0]);
  assign nor_1050_nl = ~(nor_tmp_291 | (fsm_output[8]));
  assign mux_1272_nl = MUX_s_1_2_2(mux_1271_nl, nor_1050_nl, fsm_output[5]);
  assign mux_1268_nl = MUX_s_1_2_2(and_dcpl_61, mux_528_cse, or_3185_cse);
  assign mux_1267_nl = MUX_s_1_2_2((~ (fsm_output[8])), mux_tmp_960, fsm_output[0]);
  assign mux_1269_nl = MUX_s_1_2_2((~ mux_1268_nl), mux_1267_nl, fsm_output[5]);
  assign mux_1273_nl = MUX_s_1_2_2(mux_1272_nl, mux_1269_nl, fsm_output[3]);
  assign nor_1325_nl = ~((fsm_output[6]) | mux_1273_nl);
  assign nor_1326_nl = ~((fsm_output[5]) | and_1474_cse | (fsm_output[2]) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign nor_1327_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[1])) | (fsm_output[2])
      | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1265_nl = MUX_s_1_2_2(nor_1326_nl, nor_1327_nl, fsm_output[3]);
  assign nor_1328_nl = ~(nor_1106_cse | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1329_nl = ~(and_1474_cse | (~ (fsm_output[2])) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign mux_1263_nl = MUX_s_1_2_2(nor_1328_nl, nor_1329_nl, fsm_output[5]);
  assign nor_1330_nl = ~((~(and_1572_cse | (fsm_output[4]))) | (fsm_output[8]));
  assign nor_1331_nl = ~((fsm_output[0]) | (fsm_output[1]) | (fsm_output[2]) | (~
      (fsm_output[4])) | (fsm_output[8]));
  assign mux_1262_nl = MUX_s_1_2_2(nor_1330_nl, nor_1331_nl, fsm_output[5]);
  assign mux_1264_nl = MUX_s_1_2_2(mux_1263_nl, mux_1262_nl, fsm_output[3]);
  assign mux_1266_nl = MUX_s_1_2_2(mux_1265_nl, mux_1264_nl, fsm_output[6]);
  assign GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c0 = MUX_s_1_2_2(nor_1325_nl, mux_1266_nl,
      fsm_output[7]);
  assign nor_1053_cse = ~((~ (fsm_output[6])) | (~ (fsm_output[0])) | (fsm_output[1])
      | (~ (fsm_output[2])) | (fsm_output[4]));
  assign nor_1054_nl = ~((fsm_output[6]) | (fsm_output[0]) | (~ (fsm_output[1]))
      | (fsm_output[2]) | (~ (fsm_output[4])));
  assign mux_1275_nl = MUX_s_1_2_2(nor_1053_cse, nor_1054_nl, fsm_output[7]);
  assign nor_1055_nl = ~((fsm_output[7]) | (~ (fsm_output[6])) | (~ (fsm_output[0]))
      | (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[4]));
  assign mux_1276_nl = MUX_s_1_2_2(mux_1275_nl, nor_1055_nl, CACHE_UPDATE_LOOP_1_and_tmp);
  assign GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c1 = mux_1276_nl & and_dcpl_1 & (fsm_output[3]);
  assign or_2199_nl = (~ (fsm_output[3])) | (~ (fsm_output[2])) | (fsm_output[0])
      | (~ (fsm_output[6])) | (fsm_output[7]);
  assign or_2198_nl = (fsm_output[2]) | (fsm_output[0]) | (fsm_output[6]) | (~ (fsm_output[7]));
  assign mux_1279_nl = MUX_s_1_2_2(or_2199_nl, or_2198_nl, fsm_output[5]);
  assign or_3169_nl = (fsm_output[4]) | mux_1279_nl;
  assign or_2195_nl = (~ (fsm_output[2])) | (fsm_output[0]) | (fsm_output[6]) | (~
      (fsm_output[7]));
  assign or_2193_nl = (~ CACHE_UPDATE_LOOP_1_and_tmp) | (fsm_output[0]) | (fsm_output[6])
      | (~ (fsm_output[7]));
  assign mux_1277_nl = MUX_s_1_2_2(or_2193_nl, or_2249_cse, fsm_output[2]);
  assign mux_1278_nl = MUX_s_1_2_2(or_2195_nl, mux_1277_nl, fsm_output[3]);
  assign or_3170_nl = (fsm_output[5:4]!=2'b01) | mux_1278_nl;
  assign mux_1280_nl = MUX_s_1_2_2(or_3169_nl, or_3170_nl, fsm_output[1]);
  assign GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c2 = ~(mux_1280_nl | (fsm_output[8]));
  assign GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c3 = and_dcpl_203 & and_dcpl_237;
  assign and_601_nl = (fsm_output[5]) & ((((fsm_output[1:0]!=2'b10)) & (fsm_output[2]))
      | (fsm_output[4]));
  assign mux_1283_nl = MUX_s_1_2_2(and_1762_cse, and_601_nl, fsm_output[3]);
  assign or_2203_nl = nor_593_cse | (fsm_output[4]);
  assign mux_1282_nl = MUX_s_1_2_2(mux_tmp_1281, or_2203_nl, fsm_output[0]);
  assign nor_1060_nl = ~((fsm_output[3]) | (fsm_output[5]) | mux_1282_nl);
  assign mux_1284_nl = MUX_s_1_2_2(mux_1283_nl, nor_1060_nl, fsm_output[6]);
  assign GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c6 = mux_1284_nl & and_dcpl_295;
  assign attention_abs_qr_35_0_lpi_1_dfm_mx0c1 = and_dcpl_192 & and_dcpl_564 & (~((fsm_output[7])
      | (operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1[35])));
  assign nor_1102_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (~ (fsm_output[1])) | (fsm_output[8]) | (~ (fsm_output[0])) | (fsm_output[2])
      | (~ (fsm_output[6])));
  assign nor_1099_nl = ~((fsm_output[1]) | (fsm_output[8]) | (fsm_output[0]) | (~
      (fsm_output[2])) | (fsm_output[6]));
  assign nor_1100_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[8])) | (~ LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4)
      | (fsm_output[0]) | (~ (fsm_output[2])) | (fsm_output[6]));
  assign mux_1401_nl = MUX_s_1_2_2(nor_1099_nl, nor_1100_nl, fsm_output[3]);
  assign nor_1101_nl = ~((fsm_output[3]) | (~ (fsm_output[1])) | (fsm_output[8])
      | (~ (fsm_output[0])) | (fsm_output[2]) | (~ (fsm_output[6])));
  assign mux_1402_nl = MUX_s_1_2_2(mux_1401_nl, nor_1101_nl, fsm_output[7]);
  assign and_1635_nl = (fsm_output[5]) & mux_1402_nl;
  assign RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c1 = MUX_s_1_2_2(nor_1102_nl, and_1635_nl,
      fsm_output[4]);
  assign mux_1407_nl = MUX_s_1_2_2((~ nor_tmp_285), and_1570_cse, fsm_output[5]);
  assign mux_1408_nl = MUX_s_1_2_2((~ (fsm_output[5])), mux_1407_nl, fsm_output[3]);
  assign mux_1409_nl = MUX_s_1_2_2(mux_tmp_1027, mux_1408_nl, LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4);
  assign RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c4 = (~ mux_1409_nl) & and_dcpl_413;
  assign mux_1447_nl = MUX_s_1_2_2(or_270_cse, or_255_cse, and_1474_cse);
  assign and_1642_nl = (fsm_output[6]) & (fsm_output[3]) & (~ mux_1447_nl);
  assign mux_1444_nl = MUX_s_1_2_2(and_dcpl_364, (fsm_output[4]), fsm_output[1]);
  assign mux_1445_nl = MUX_s_1_2_2((~ mux_1444_nl), or_tmp_1221, fsm_output[0]);
  assign mux_1442_nl = MUX_s_1_2_2(or_tmp_11, mux_tmp_87, fsm_output[1]);
  assign mux_1443_nl = MUX_s_1_2_2(mux_1442_nl, mux_tmp_834, fsm_output[0]);
  assign mux_1446_nl = MUX_s_1_2_2(mux_1445_nl, mux_1443_nl, fsm_output[3]);
  assign nor_1111_nl = ~((fsm_output[6]) | mux_1446_nl);
  assign mux_1448_nl = MUX_s_1_2_2(and_1642_nl, nor_1111_nl, fsm_output[7]);
  assign CACHE_UPDATE_LOOP_3_k_2_0_sva_1_mx0c1 = mux_1448_nl & and_dcpl_1;
  assign nor_1118_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[0])) | (~ (fsm_output[6]))
      | (fsm_output[5]) | (fsm_output[8]));
  assign nor_1119_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[0])) | (fsm_output[6])
      | (fsm_output[5]) | (~ (fsm_output[8])));
  assign mux_1464_nl = MUX_s_1_2_2(nor_1118_nl, nor_1119_nl, fsm_output[4]);
  assign and_1644_nl = (~((fsm_output[1]) | (~ (fsm_output[3])))) & mux_1464_nl;
  assign nor_1120_nl = ~((~ (fsm_output[3])) | (fsm_output[4]) | (fsm_output[2])
      | (fsm_output[0]) | (fsm_output[6]) | (~ (fsm_output[5])) | (fsm_output[8]));
  assign or_2363_nl = (z_out_5[2]) | (~ (fsm_output[0])) | (~ (fsm_output[6])) |
      (fsm_output[5]) | (fsm_output[8]);
  assign or_2362_nl = (z_out_5[2]) | (fsm_output[0]) | (fsm_output[6]) | (~ (fsm_output[5]))
      | (fsm_output[8]);
  assign mux_1461_nl = MUX_s_1_2_2(or_2363_nl, or_2362_nl, fsm_output[2]);
  assign nor_1121_nl = ~((fsm_output[4]) | mux_1461_nl);
  assign nor_1122_nl = ~((fsm_output[0]) | (~ (fsm_output[6])) | (fsm_output[5])
      | (fsm_output[8]));
  assign nor_1123_nl = ~((~ (fsm_output[0])) | (fsm_output[6]) | (fsm_output[5])
      | (fsm_output[8]));
  assign mux_1459_nl = MUX_s_1_2_2(nor_1122_nl, nor_1123_nl, fsm_output[2]);
  assign nor_1124_nl = ~((fsm_output[0]) | CACHE_UPDATE_LOOP_1_and_tmp | (fsm_output[6])
      | (fsm_output[5]) | (fsm_output[8]));
  assign nor_1125_nl = ~((z_out_5[2]) | (~ (fsm_output[0])) | (fsm_output[6]) | (fsm_output[5])
      | (fsm_output[8]));
  assign mux_1458_nl = MUX_s_1_2_2(nor_1124_nl, nor_1125_nl, fsm_output[2]);
  assign mux_1460_nl = MUX_s_1_2_2(mux_1459_nl, mux_1458_nl, fsm_output[4]);
  assign mux_1462_nl = MUX_s_1_2_2(nor_1121_nl, mux_1460_nl, fsm_output[3]);
  assign mux_1463_nl = MUX_s_1_2_2(nor_1120_nl, mux_1462_nl, fsm_output[1]);
  assign GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c1 = MUX_s_1_2_2(and_1644_nl, mux_1463_nl,
      fsm_output[7]);
  assign nor_1129_nl = ~((fsm_output[1]) | RESHAPE_2D_TO_3D_LOOP_2_2_and_cse | (fsm_output[8:4]!=5'b01001));
  assign nor_1130_nl = ~((~ (fsm_output[1])) | (~ (z_out_5[2])) | (fsm_output[8:4]!=5'b01100));
  assign mux_1473_nl = MUX_s_1_2_2(nor_1129_nl, nor_1130_nl, fsm_output[0]);
  assign nor_1126_nl = ~((fsm_output[8:4]!=5'b01001));
  assign nor_1127_nl = ~((~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign nor_1128_nl = ~((~ (fsm_output[7])) | (fsm_output[6]) | (fsm_output[4])
      | (fsm_output[8]));
  assign mux_1471_nl = MUX_s_1_2_2(nor_1127_nl, nor_1128_nl, fsm_output[5]);
  assign mux_1472_nl = MUX_s_1_2_2(nor_1126_nl, mux_1471_nl, z_out_5[2]);
  assign and_1646_nl = nor_366_cse & mux_1472_nl;
  assign mux_1474_nl = MUX_s_1_2_2(mux_1473_nl, and_1646_nl, fsm_output[2]);
  assign nor_1131_nl = ~((~ (fsm_output[1])) | (~ CACHE_UPDATE_LOOP_1_and_tmp) |
      (fsm_output[8:4]!=5'b01001));
  assign nor_1132_nl = ~((fsm_output[1]) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[6]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1469_nl = MUX_s_1_2_2(nor_1131_nl, nor_1132_nl, fsm_output[0]);
  assign nor_1133_nl = ~((fsm_output[5]) | (fsm_output[7]) | mux_1309_cse);
  assign nor_1134_nl = ~((fsm_output[8:4]!=5'b01000));
  assign mux_1467_nl = MUX_s_1_2_2(nor_1133_nl, nor_1134_nl, fsm_output[1]);
  assign nor_1135_nl = ~((~ (fsm_output[1])) | (~ (z_out_5[2])) | (fsm_output[8:4]!=5'b01001));
  assign mux_1468_nl = MUX_s_1_2_2(mux_1467_nl, nor_1135_nl, fsm_output[0]);
  assign mux_1470_nl = MUX_s_1_2_2(mux_1469_nl, mux_1468_nl, fsm_output[2]);
  assign GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c2 = MUX_s_1_2_2(mux_1474_nl, mux_1470_nl,
      fsm_output[3]);
  assign or_2499_nl = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b10)
      | (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd) | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  assign mux_1586_nl = MUX_s_1_2_2(nor_1026_cse, mux_tmp_1578, or_2499_nl);
  assign attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16_mx0c1 = mux_1586_nl &
      (~ (fsm_output[8])) & and_dcpl_814;
  assign nand_359_nl = ~((reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2==2'b11)
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1));
  assign mux_1592_nl = MUX_s_1_2_2(nor_1026_cse, mux_tmp_1578, nand_359_nl);
  assign attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16_mx0c1 = mux_1592_nl &
      (~ (fsm_output[8])) & and_dcpl_814;
  assign and_1811_cse = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  assign mux_2262_nl = MUX_s_1_2_2(mux_tmp_1578, (~ or_tmp_1354), and_1811_cse);
  assign mux_1594_nl = MUX_s_1_2_2(mux_2262_nl, mux_tmp_1578, or_dcpl_332);
  assign attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16_mx0c1 = mux_1594_nl &
      (~ (fsm_output[8])) & and_dcpl_814;
  assign mux_1593_nl = MUX_s_1_2_2(mux_tmp_1578, (~ or_tmp_1354), and_1811_cse);
  assign mux_1595_nl = MUX_s_1_2_2(mux_1593_nl, mux_tmp_1578, or_dcpl_342);
  assign attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16_mx0c1 = mux_1595_nl &
      (~ (fsm_output[8])) & and_dcpl_814;
  assign mux_1596_nl = MUX_s_1_2_2(nor_1026_cse, mux_tmp_1578, or_2739_cse);
  assign attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16_mx0c1 = mux_1596_nl &
      (~ (fsm_output[8])) & and_dcpl_814;
  assign and_1659_nl = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[1])
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  assign mux_1597_nl = MUX_s_1_2_2(mux_tmp_1578, (~ or_tmp_1354), and_1659_nl);
  assign mux_1598_nl = MUX_s_1_2_2(mux_1597_nl, mux_tmp_1578, reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]);
  assign attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16_mx0c1 = mux_1598_nl &
      (~ (fsm_output[8])) & and_dcpl_814;
  assign mux_1599_nl = MUX_s_1_2_2(nor_1026_cse, mux_tmp_1578, or_3039_cse);
  assign attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16_mx0c1 = mux_1599_nl &
      (~ (fsm_output[8])) & and_dcpl_814;
  assign nand_361_nl = ~(RESHAPE_2D_TO_3D_LOOP_2_2_and_cse & (fsm_output[4]) & (~
      (fsm_output[0])) & (fsm_output[7]));
  assign nand_362_nl = ~((fsm_output[4]) & (fsm_output[0]) & (fsm_output[7]));
  assign mux_1605_nl = MUX_s_1_2_2(nand_361_nl, nand_362_nl, fsm_output[3]);
  assign nor_1160_nl = ~((fsm_output[2]) | mux_1605_nl);
  assign nor_1161_nl = ~((~((fsm_output[3]) | RESHAPE_2D_TO_3D_LOOP_2_2_and_cse))
      | (~ (fsm_output[4])) | (fsm_output[0]) | (~ (fsm_output[7])));
  assign nor_1162_nl = ~((~ (fsm_output[4])) | (fsm_output[0]) | (~ (fsm_output[7])));
  assign nor_1163_nl = ~((fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[7])));
  assign mux_1603_nl = MUX_s_1_2_2(nor_1162_nl, nor_1163_nl, fsm_output[3]);
  assign mux_1604_nl = MUX_s_1_2_2(nor_1161_nl, mux_1603_nl, fsm_output[2]);
  assign mux_1606_nl = MUX_s_1_2_2(nor_1160_nl, mux_1604_nl, fsm_output[1]);
  assign nor_1164_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[7])));
  assign mux_1601_nl = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[0]);
  assign nor_1165_nl = ~((fsm_output[4:2]!=3'b010) | mux_1601_nl);
  assign mux_1602_nl = MUX_s_1_2_2(nor_1164_nl, nor_1165_nl, fsm_output[1]);
  assign mux_1607_nl = MUX_s_1_2_2(mux_1606_nl, mux_1602_nl, fsm_output[6]);
  assign APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c0 = mux_1607_nl & and_dcpl_1;
  assign mux_1608_nl = MUX_s_1_2_2(and_1555_cse, nor_749_cse, fsm_output[3]);
  assign APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c2 = mux_1608_nl & and_dcpl_201
      & and_dcpl_577 & and_dcpl_45;
  assign and_1666_nl = (fsm_output[4]) & (~(nor_1106_cse | (~ (fsm_output[3])) |
      (fsm_output[6])));
  assign nor_1169_nl = ~(((fsm_output[4:0]==5'b11111)) | (fsm_output[6]));
  assign mux_1610_nl = MUX_s_1_2_2(and_1666_nl, nor_1169_nl, fsm_output[5]);
  assign and_1667_nl = (fsm_output[8]) & mux_1610_nl;
  assign nor_1170_nl = ~((~ (fsm_output[1])) | (fsm_output[2]) | (~ (fsm_output[3]))
      | (fsm_output[6]));
  assign nor_1171_nl = ~((fsm_output[0]) | (fsm_output[1]) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (~ (fsm_output[6])));
  assign mux_1609_nl = MUX_s_1_2_2(nor_1170_nl, nor_1171_nl, fsm_output[4]);
  assign and_1668_nl = (~((fsm_output[8]) | (~ (fsm_output[5])))) & mux_1609_nl;
  assign APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c3 = MUX_s_1_2_2(and_1667_nl,
      and_1668_nl, fsm_output[7]);
  assign or_2541_nl = (fsm_output[3]) | (fsm_output[0]) | (~ (fsm_output[4]));
  assign mux_1614_nl = MUX_s_1_2_2(or_2541_nl, or_tmp_1392, fsm_output[6]);
  assign or_3189_nl = or_tmp_1392 | (~ (fsm_output[6]));
  assign mux_1615_nl = MUX_s_1_2_2(mux_1614_nl, or_3189_nl, RESHAPE_2D_TO_3D_LOOP_2_2_and_cse);
  assign APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c4 = (~ mux_1615_nl) & and_dcpl_226
      & and_dcpl_885;
  assign apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c1 = and_dcpl_732
      & and_dcpl_604;
  assign apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c8 = and_dcpl_743
      & and_dcpl_551 & and_dcpl_728;
  assign apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1 = and_dcpl_732
      & and_dcpl_1000;
  assign attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c1 = and_dcpl_732 & and_dcpl_721;
  assign attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c6 = and_dcpl_743 & and_dcpl_552;
  assign attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0_mx0c1 = and_dcpl_732 & and_dcpl_591
      & and_dcpl_462;
  assign or_2762_nl = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b11)
      | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  assign mux_2060_nl = MUX_s_1_2_2(nor_1026_cse, mux_tmp_1578, or_2762_nl);
  assign apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16_mx0c1 = mux_2060_nl
      & (~ (fsm_output[8])) & and_dcpl_814;
  assign or_2768_nl = (~ reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd!=3'b001);
  assign mux_2069_nl = MUX_s_1_2_2(or_1983_cse, mux_tmp_1562, or_2768_nl);
  assign apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16_mx0c1 = (~(mux_2069_nl
      | (fsm_output[8]))) & and_dcpl_748;
  assign and_1781_cse = (fsm_output[8]) & (~(and_1782_cse | (fsm_output[6:5]!=2'b00)));
  assign and_1778_nl = (((fsm_output[1:0]==2'b11) & (z_out_5[2])) | (fsm_output[5]))
      & (fsm_output[6]);
  assign mux_2138_nl = MUX_s_1_2_2(and_1778_nl, (fsm_output[6]), fsm_output[2]);
  assign or_1238_nl = (fsm_output[6:5]!=2'b00);
  assign mux_2136_nl = MUX_s_1_2_2(or_1238_nl, (fsm_output[5]), or_3163_cse);
  assign mux_2137_nl = MUX_s_1_2_2((fsm_output[6]), mux_2136_nl, nor_593_cse);
  assign mux_2139_cse = MUX_s_1_2_2(mux_2138_nl, mux_2137_nl, fsm_output[3]);
  assign or_2858_cse = nor_305_cse | (fsm_output[6]);
  assign or_2856_cse = nor_1026_cse | (fsm_output[6]);
  assign and_1780_nl = (~(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 & (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0])
      & (fsm_output[0]) & (fsm_output[5]))) & (fsm_output[6]);
  assign mux_2132_nl = MUX_s_1_2_2(and_1780_nl, (fsm_output[6]), or_dcpl_672);
  assign mux_2133_nl = MUX_s_1_2_2(or_2856_cse, mux_2132_nl, fsm_output[1]);
  assign mux_2134_nl = MUX_s_1_2_2(or_2858_cse, mux_2133_nl, fsm_output[2]);
  assign mux_2135_nl = MUX_s_1_2_2(mux_2134_nl, (fsm_output[6]), fsm_output[3]);
  assign mux_2140_nl = MUX_s_1_2_2(mux_2139_cse, mux_2135_nl, fsm_output[4]);
  assign nor_1234_nl = ~((fsm_output[8]) | (~ mux_2140_nl));
  assign attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c1 = MUX_s_1_2_2(and_1781_cse,
      nor_1234_nl, fsm_output[7]);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c9 = and_dcpl_360 &
      and_dcpl_355 & and_dcpl_539;
  assign attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx0c7 = and_dcpl_360 &
      and_dcpl_355 & and_dcpl_651;
  assign attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx0c7 = and_dcpl_360 &
      and_dcpl_355 & and_dcpl_656;
  assign and_1790_cse = (~((fsm_output[0]) & (fsm_output[5]))) & (fsm_output[6]);
  assign mux_2183_nl = MUX_s_1_2_2(and_1790_cse, (fsm_output[6]), or_2671_cse);
  assign mux_2184_nl = MUX_s_1_2_2(or_2856_cse, mux_2183_nl, fsm_output[1]);
  assign mux_2185_nl = MUX_s_1_2_2(or_2858_cse, mux_2184_nl, fsm_output[2]);
  assign mux_2186_nl = MUX_s_1_2_2(mux_2185_nl, (fsm_output[6]), fsm_output[3]);
  assign mux_2191_nl = MUX_s_1_2_2(mux_2139_cse, mux_2186_nl, fsm_output[4]);
  assign nor_1261_nl = ~((fsm_output[8]) | (~ mux_2191_nl));
  assign attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c1 = MUX_s_1_2_2(and_1781_cse,
      nor_1261_nl, fsm_output[7]);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c9 = and_dcpl_360 &
      and_dcpl_513 & and_dcpl_354;
  assign attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx0c7 = and_dcpl_360 &
      and_dcpl_513 & and_dcpl_458;
  assign attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx0c7 = and_dcpl_360 &
      and_dcpl_513 & and_dcpl_651;
  assign attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx0c7 = and_dcpl_360 &
      and_dcpl_513 & and_dcpl_656;
  assign mux_2211_nl = MUX_s_1_2_2(and_1790_cse, (fsm_output[6]), or_2486_cse);
  assign mux_2212_nl = MUX_s_1_2_2(or_2856_cse, mux_2211_nl, fsm_output[1]);
  assign mux_2213_nl = MUX_s_1_2_2(or_2858_cse, mux_2212_nl, fsm_output[2]);
  assign mux_2214_nl = MUX_s_1_2_2(mux_2213_nl, (fsm_output[6]), fsm_output[3]);
  assign mux_2219_nl = MUX_s_1_2_2(mux_2139_cse, mux_2214_nl, fsm_output[4]);
  assign nor_1299_nl = ~((fsm_output[8]) | (~ mux_2219_nl));
  assign attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c1 = MUX_s_1_2_2(and_1781_cse,
      nor_1299_nl, fsm_output[7]);
  assign attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c9 = and_dcpl_360 &
      and_dcpl_355 & and_dcpl_512;
  assign attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx0c7 = and_dcpl_360 &
      and_dcpl_355 & and_dcpl_525;
  assign attention_abs_4_qr_35_0_lpi_1_dfm_mx0c1 = and_dcpl_362 & and_dcpl_198 &
      (fsm_output[7:6]==2'b11) & (~ (operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1[35]));
  assign GEMM_3D_FLOAT_LOOP_4_l_and_ssc = attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1
      & (GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c0 | GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c1
      | GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c2 | GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c3
      | and_dcpl_193 | and_dcpl_349 | GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c6);
  assign GEMM_3D_FLOAT_LOOP_4_l_or_2_cse = GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c1
      | and_dcpl_349;
  assign CACHE_UPDATE_LOOP_3_mux_3_nl = MUX_v_40_16_2(attention_2_1_16_16_4_4_k_embed_0_0_0_sva_1,
      attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1, attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1,
      attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1, attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1,
      attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1, attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1,
      attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1,
      attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1,
      attention_2_1_16_16_4_4_k_embed_2_0_3_sva_1, attention_2_1_16_16_4_4_k_embed_3_0_0_sva_1,
      attention_2_1_16_16_4_4_k_embed_3_0_1_sva_1, attention_2_1_16_16_4_4_k_embed_3_0_2_sva_1,
      attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1, {reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1});
  assign and_369_nl = and_dcpl_322 & and_dcpl_319 & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2==2'b10);
  assign attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d = MUX_v_40_2_2(({{21{CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_itm[18]}},
      CACHE_UPDATE_LOOP_3_qif_read_rom_k_cache_rom_map_1_itm}), CACHE_UPDATE_LOOP_3_mux_3_nl,
      and_369_nl);
  assign nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_nl = conv_u2u_2_3(TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_sdt_1[2:1])
      + conv_u2u_2_3({reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_nl = nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_nl[2:0];
  assign attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d = {TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_nl
      , (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_sdt_1[0]) , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1};
  assign attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_pff = and_dcpl_328;
  assign nl_CACHE_UPDATE_LOOP_3_acc_nl = conv_u2u_2_3(CACHE_UPDATE_LOOP_3_acc_sdt_1[2:1])
      + conv_u2u_2_3({reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign CACHE_UPDATE_LOOP_3_acc_nl = nl_CACHE_UPDATE_LOOP_3_acc_nl[2:0];
  assign attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d = {CACHE_UPDATE_LOOP_3_acc_nl
      , (CACHE_UPDATE_LOOP_3_acc_sdt_1[0]) , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0
      , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1};
  assign attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_pff = and_dcpl_318;
  assign CACHE_UPDATE_LOOP_3_1_mux_2_nl = MUX_v_24_16_2(attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16, {reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign CACHE_UPDATE_LOOP_3_1_CACHE_UPDATE_LOOP_3_1_mux_nl = MUX_v_24_2_2((signext_24_4(CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_sdt[19:16])),
      CACHE_UPDATE_LOOP_3_1_mux_2_nl, and_362_ssc);
  assign CACHE_UPDATE_LOOP_3_1_mux_3_nl = MUX_v_16_16_2(attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0, {reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign CACHE_UPDATE_LOOP_3_1_CACHE_UPDATE_LOOP_3_1_mux_1_nl = MUX_v_16_2_2((CACHE_UPDATE_LOOP_3_1_qif_read_rom_v_cache_rom_map_1_sdt[15:0]),
      CACHE_UPDATE_LOOP_3_1_mux_3_nl, and_362_ssc);
  assign attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d = {CACHE_UPDATE_LOOP_3_1_CACHE_UPDATE_LOOP_3_1_mux_nl
      , CACHE_UPDATE_LOOP_3_1_CACHE_UPDATE_LOOP_3_1_mux_1_nl};
  assign nl_GEMM_3D_FLOAT_LOOP_4_1_acc_13_nl = conv_u2u_2_3(GEMM_3D_FLOAT_LOOP_4_1_acc_12_sdt_1[2:1])
      + conv_u2u_2_3({reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign GEMM_3D_FLOAT_LOOP_4_1_acc_13_nl = nl_GEMM_3D_FLOAT_LOOP_4_1_acc_13_nl[2:0];
  assign attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d = {GEMM_3D_FLOAT_LOOP_4_1_acc_13_nl
      , (GEMM_3D_FLOAT_LOOP_4_1_acc_12_sdt_1[0]) , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1};
  assign attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_pff = and_dcpl_316;
  assign attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d = {GEMM_3D_FLOAT_LOOP_3_acc_6_tmp
      , (z_out_11[0]) , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1};
  assign nl_GEMM_3D_FLOAT_LOOP_4_acc_nl = conv_u2u_2_3(GEMM_3D_FLOAT_LOOP_4_acc_sdt_1[2:1])
      + conv_u2u_2_3({reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign GEMM_3D_FLOAT_LOOP_4_acc_nl = nl_GEMM_3D_FLOAT_LOOP_4_acc_nl[2:0];
  assign attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d = {GEMM_3D_FLOAT_LOOP_4_acc_nl
      , (GEMM_3D_FLOAT_LOOP_4_acc_sdt_1[0]) , (GEMM_3D_FLOAT_LOOP_4_acc_13_sdt_1[0])
      , (z_out_11[0])};
  assign attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_pff = and_dcpl_313;
  assign attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d = {TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_16_psp_1
      , (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]) , reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2};
  assign attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_pff = and_dcpl_289 &
      and_dcpl_237;
  assign and_dcpl_1233 = and_dcpl_222 & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd;
  assign and_dcpl_1248 = (fsm_output[4:0]==5'b01111) & and_dcpl_1 & (fsm_output[7:6]==2'b10);
  assign and_dcpl_1261 = and_dcpl_61 & (fsm_output[2]) & (fsm_output[1]) & (fsm_output[0])
      & (fsm_output[3]) & (~ (fsm_output[5])) & (~ (fsm_output[6])) & (fsm_output[7]);
  assign nor_1345_nl = ~((fsm_output[6]) | (fsm_output[2]) | or_dcpl_959);
  assign nor_1346_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[2])) | (fsm_output[4])
      | (fsm_output[8]));
  assign mux_2299_nl = MUX_s_1_2_2(nor_1345_nl, nor_1346_nl, fsm_output[7]);
  assign and_dcpl_1273 = mux_2299_nl & (~ (fsm_output[1])) & (fsm_output[0]) & (fsm_output[3])
      & (~ (fsm_output[5]));
  assign and_dcpl_1294 = nor_1314_cse & (~ (fsm_output[1])) & (fsm_output[0]) & (~
      (fsm_output[5])) & (fsm_output[7]);
  assign and_dcpl_1363 = (fsm_output==9'b011110101);
  assign and_dcpl_1371 = (~ (fsm_output[8])) & (fsm_output[4]) & (~ (fsm_output[1]))
      & (fsm_output[2]) & (~ (fsm_output[0])) & and_dcpl_198 & (fsm_output[7:6]==2'b10);
  assign and_dcpl_1379 = and_dcpl_61 & (fsm_output[1]) & and_1555_cse & and_dcpl_181
      & (fsm_output[7:6]==2'b01);
  assign and_dcpl_1385 = (fsm_output[8]) & (fsm_output[4]) & (fsm_output[1]) & and_1555_cse
      & and_dcpl_181 & nor_973_cse;
  assign and_dcpl_1391 = and_dcpl_61 & (fsm_output[1]);
  assign and_dcpl_1392 = and_dcpl_1391 & nor_749_cse;
  assign and_dcpl_1393 = and_dcpl_1392 & and_dcpl_209;
  assign and_dcpl_1396 = and_dcpl_201 & (fsm_output[1]);
  assign and_dcpl_1398 = and_dcpl_1396 & (~ (fsm_output[2])) & (fsm_output[0]) &
      and_dcpl_209;
  assign and_dcpl_1401 = (fsm_output[2]) & (~ (fsm_output[0]));
  assign and_dcpl_1403 = and_dcpl_1396 & and_dcpl_1401 & (~ (fsm_output[3])) & (fsm_output[5])
      & nor_973_cse;
  assign and_dcpl_1406 = and_dcpl_181 & (fsm_output[7:6]==2'b01);
  assign and_dcpl_1407 = and_dcpl_1392 & and_dcpl_1406;
  assign and_dcpl_1410 = and_dcpl_1391 & and_1555_cse & and_dcpl_1406;
  assign and_dcpl_1415 = and_dcpl_201 & (~ (fsm_output[1])) & and_dcpl_1401 & and_dcpl_198
      & and_dcpl_45;
  assign nor_1378_nl = ~((~ (fsm_output[5])) | (fsm_output[2]));
  assign nor_1379_nl = ~((fsm_output[5]) | (~ (fsm_output[2])));
  assign mux_2288_nl = MUX_s_1_2_2(nor_1378_nl, nor_1379_nl, fsm_output[6]);
  assign and_dcpl_1420 = mux_2288_nl & and_dcpl_61 & (fsm_output[1]) & (fsm_output[0])
      & (~ (fsm_output[3])) & (fsm_output[7]);
  assign and_dcpl_1425 = and_dcpl_61 & (~ (fsm_output[1])) & and_1555_cse & (fsm_output[3])
      & (fsm_output[5]) & and_dcpl_45;
  assign and_dcpl_1427 = and_dcpl_181 & (fsm_output[7:6]==2'b11);
  assign and_dcpl_1429 = and_dcpl_1391 & and_dcpl_1401 & and_dcpl_1427;
  assign and_dcpl_1431 = and_dcpl_1396 & and_1555_cse & and_dcpl_1427;
  assign and_dcpl_1436 = (fsm_output[8]) & (fsm_output[4]) & (fsm_output[1]) & nor_749_cse
      & and_dcpl_181 & nor_973_cse;
  assign RMS_NORM_LOOP_1_1_or_3_ssc = and_dcpl_1403 | and_dcpl_1410 | and_dcpl_1420
      | and_dcpl_1425 | and_dcpl_1429;
  assign RMS_NORM_LOOP_1_1_or_1_ssc = and_dcpl_1407 | and_dcpl_1436;
  assign or_3261_nl = (fsm_output[3]) | nand_240_cse;
  assign or_3235_nl = (fsm_output[2]) | (fsm_output[1]) | (fsm_output[4]);
  assign mux_2290_nl = MUX_s_1_2_2(or_3235_nl, or_tmp_1128, fsm_output[0]);
  assign mux_2291_nl = MUX_s_1_2_2(mux_2290_nl, mux_1513_cse, fsm_output[3]);
  assign mux_2292_nl = MUX_s_1_2_2(or_3261_nl, mux_2291_nl, fsm_output[5]);
  assign and_dcpl_1447 = (~ mux_2292_nl) & and_dcpl_307 & (fsm_output[7]);
  assign RMS_NORM_LOOP_1_1_or_2_ssc = and_dcpl_1407 | and_dcpl_1425 | and_dcpl_1429;
  assign and_1908_cse = and_dcpl_61 & (fsm_output[1]) & (fsm_output[2]) & (~ (fsm_output[0]))
      & (fsm_output[3]) & (~ (fsm_output[5])) & (fsm_output[6]) & (~ (fsm_output[7]));
  assign mux_2266_nl = MUX_s_1_2_2(nor_176_cse, and_1651_cse, fsm_output[2]);
  assign nor_1348_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[1])) | (fsm_output[4]));
  assign mux_2267_nl = MUX_s_1_2_2(mux_2266_nl, nor_1348_nl, fsm_output[3]);
  assign CACHE_UPDATE_LOOP_3_or_cse = (mux_2267_nl & (~ (fsm_output[8])) & (fsm_output[0])
      & (~ (fsm_output[5])) & and_dcpl_45) | and_1908_cse;
  assign nor_1350_nl = ~((fsm_output[6]) | (fsm_output[0]) | (fsm_output[2]) | (~
      and_1651_cse));
  assign mux_2268_nl = MUX_s_1_2_2(nor_1053_cse, nor_1350_nl, fsm_output[7]);
  assign nand_394_nl = ~((fsm_output[3]) & (fsm_output[1]) & (fsm_output[4]));
  assign mux_2270_nl = MUX_s_1_2_2(nand_394_nl, or_tmp_704, fsm_output[5]);
  assign CACHE_UPDATE_LOOP_3_or_1_cse = (mux_2268_nl & (~ (fsm_output[8])) & (fsm_output[3])
      & (~ (fsm_output[5]))) | ((~(mux_2270_nl | (fsm_output[8]))) & (~ (fsm_output[2]))
      & (fsm_output[0]) & and_dcpl_45);
  assign RMS_NORM_LOOP_1_1_or_5_cse = and_dcpl_1398 | and_dcpl_1403 | and_dcpl_1431;
  assign RMS_NORM_LOOP_1_1_nor_seb = ~(and_dcpl_1398 | and_dcpl_1431);
  assign RMS_NORM_LOOP_1_1_or_4_itm = and_dcpl_1398 | and_dcpl_1431;
  assign nand_398_nl = ~((fsm_output[1]) & (fsm_output[4]));
  assign mux_2286_nl = MUX_s_1_2_2(or_tmp_11, nand_398_nl, fsm_output[0]);
  assign nor_1368_nl = ~((fsm_output[3]) | mux_2286_nl);
  assign nor_1369_nl = ~((fsm_output[4:0]!=5'b01011));
  assign mux_2287_nl = MUX_s_1_2_2(nor_1368_nl, nor_1369_nl, fsm_output[6]);
  assign GEMM_3D_FLOAT_LOOP_1_or_ssc = and_1908_cse | (mux_2287_nl & and_dcpl_1 &
      (fsm_output[7]));
  always @(posedge clk) begin
    if ( rst ) begin
      strm_out_rsci_idat_17_10 <= 8'b00000000;
      strm_out_rsci_idat_9 <= 1'b0;
      strm_out_rsci_idat_8 <= 1'b0;
      strm_out_rsci_idat_7 <= 1'b0;
      strm_out_rsci_idat_6 <= 1'b0;
      strm_out_rsci_idat_5 <= 1'b0;
      strm_out_rsci_idat_4 <= 1'b0;
      strm_out_rsci_idat_3 <= 1'b0;
      strm_out_rsci_idat_2 <= 1'b0;
      strm_out_rsci_idat_31_18 <= 14'b00000000000000;
    end
    else if ( for_1_for_and_cse ) begin
      strm_out_rsci_idat_17_10 <= MUX_v_8_16_2((output_0_0_sva_2_15_0[15:8]), output_0_1_sva_2_15_8,
          (output_0_2_sva_2_15_0[15:8]), (output_0_3_sva_2_15_0[15:8]), (output_0_4_sva_2_15_0[15:8]),
          (output_0_5_sva_2_15_0[15:8]), (output_0_6_sva_2_15_0[15:8]), (output_0_7_sva_2_15_0[15:8]),
          (output_0_8_sva_2_15_0[15:8]), (output_0_9_sva_2_15_0[15:8]), (output_0_10_sva_2_15_0[15:8]),
          (output_0_11_sva_2_15_0[15:8]), (output_0_12_sva_2_15_0[15:8]), (output_0_13_sva_2_15_0[15:8]),
          (output_0_14_sva_2_15_0[15:8]), (output_0_15_sva_2_15_0[15:8]), {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
          , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
      strm_out_rsci_idat_9 <= MUX_s_1_16_2((output_0_0_sva_2_15_0[7]), output_0_1_sva_2_7,
          (output_0_2_sva_2_15_0[7]), (output_0_3_sva_2_15_0[7]), (output_0_4_sva_2_15_0[7]),
          (output_0_5_sva_2_15_0[7]), (output_0_6_sva_2_15_0[7]), (output_0_7_sva_2_15_0[7]),
          (output_0_8_sva_2_15_0[7]), (output_0_9_sva_2_15_0[7]), (output_0_10_sva_2_15_0[7]),
          (output_0_11_sva_2_15_0[7]), (output_0_12_sva_2_15_0[7]), (output_0_13_sva_2_15_0[7]),
          (output_0_14_sva_2_15_0[7]), (output_0_15_sva_2_15_0[7]), {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
          , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
      strm_out_rsci_idat_8 <= MUX_s_1_16_2((output_0_0_sva_2_15_0[6]), output_0_1_sva_2_6,
          (output_0_2_sva_2_15_0[6]), (output_0_3_sva_2_15_0[6]), (output_0_4_sva_2_15_0[6]),
          (output_0_5_sva_2_15_0[6]), (output_0_6_sva_2_15_0[6]), (output_0_7_sva_2_15_0[6]),
          (output_0_8_sva_2_15_0[6]), (output_0_9_sva_2_15_0[6]), (output_0_10_sva_2_15_0[6]),
          (output_0_11_sva_2_15_0[6]), (output_0_12_sva_2_15_0[6]), (output_0_13_sva_2_15_0[6]),
          (output_0_14_sva_2_15_0[6]), (output_0_15_sva_2_15_0[6]), {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
          , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
      strm_out_rsci_idat_7 <= MUX_s_1_16_2((output_0_0_sva_2_15_0[5]), output_0_1_sva_2_5,
          (output_0_2_sva_2_15_0[5]), (output_0_3_sva_2_15_0[5]), (output_0_4_sva_2_15_0[5]),
          (output_0_5_sva_2_15_0[5]), (output_0_6_sva_2_15_0[5]), (output_0_7_sva_2_15_0[5]),
          (output_0_8_sva_2_15_0[5]), (output_0_9_sva_2_15_0[5]), (output_0_10_sva_2_15_0[5]),
          (output_0_11_sva_2_15_0[5]), (output_0_12_sva_2_15_0[5]), (output_0_13_sva_2_15_0[5]),
          (output_0_14_sva_2_15_0[5]), (output_0_15_sva_2_15_0[5]), {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
          , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
      strm_out_rsci_idat_6 <= MUX_s_1_16_2((output_0_0_sva_2_15_0[4]), output_0_1_sva_2_4,
          (output_0_2_sva_2_15_0[4]), (output_0_3_sva_2_15_0[4]), (output_0_4_sva_2_15_0[4]),
          (output_0_5_sva_2_15_0[4]), (output_0_6_sva_2_15_0[4]), (output_0_7_sva_2_15_0[4]),
          (output_0_8_sva_2_15_0[4]), (output_0_9_sva_2_15_0[4]), (output_0_10_sva_2_15_0[4]),
          (output_0_11_sva_2_15_0[4]), (output_0_12_sva_2_15_0[4]), (output_0_13_sva_2_15_0[4]),
          (output_0_14_sva_2_15_0[4]), (output_0_15_sva_2_15_0[4]), {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
          , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
      strm_out_rsci_idat_5 <= MUX_s_1_16_2((output_0_0_sva_2_15_0[3]), output_0_1_sva_2_3,
          (output_0_2_sva_2_15_0[3]), (output_0_3_sva_2_15_0[3]), (output_0_4_sva_2_15_0[3]),
          (output_0_5_sva_2_15_0[3]), (output_0_6_sva_2_15_0[3]), (output_0_7_sva_2_15_0[3]),
          (output_0_8_sva_2_15_0[3]), (output_0_9_sva_2_15_0[3]), (output_0_10_sva_2_15_0[3]),
          (output_0_11_sva_2_15_0[3]), (output_0_12_sva_2_15_0[3]), (output_0_13_sva_2_15_0[3]),
          (output_0_14_sva_2_15_0[3]), (output_0_15_sva_2_15_0[3]), {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
          , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
      strm_out_rsci_idat_4 <= MUX_s_1_16_2((output_0_0_sva_2_15_0[2]), output_0_1_sva_2_2,
          (output_0_2_sva_2_15_0[2]), (output_0_3_sva_2_15_0[2]), (output_0_4_sva_2_15_0[2]),
          (output_0_5_sva_2_15_0[2]), (output_0_6_sva_2_15_0[2]), (output_0_7_sva_2_15_0[2]),
          (output_0_8_sva_2_15_0[2]), (output_0_9_sva_2_15_0[2]), (output_0_10_sva_2_15_0[2]),
          (output_0_11_sva_2_15_0[2]), (output_0_12_sva_2_15_0[2]), (output_0_13_sva_2_15_0[2]),
          (output_0_14_sva_2_15_0[2]), (output_0_15_sva_2_15_0[2]), {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
          , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
      strm_out_rsci_idat_3 <= MUX_s_1_16_2((output_0_0_sva_2_15_0[1]), output_0_1_sva_2_1,
          (output_0_2_sva_2_15_0[1]), (output_0_3_sva_2_15_0[1]), (output_0_4_sva_2_15_0[1]),
          (output_0_5_sva_2_15_0[1]), (output_0_6_sva_2_15_0[1]), (output_0_7_sva_2_15_0[1]),
          (output_0_8_sva_2_15_0[1]), (output_0_9_sva_2_15_0[1]), (output_0_10_sva_2_15_0[1]),
          (output_0_11_sva_2_15_0[1]), (output_0_12_sva_2_15_0[1]), (output_0_13_sva_2_15_0[1]),
          (output_0_14_sva_2_15_0[1]), (output_0_15_sva_2_15_0[1]), {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
          , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
      strm_out_rsci_idat_2 <= MUX_s_1_16_2((output_0_0_sva_2_15_0[0]), output_0_1_sva_2_0,
          (output_0_2_sva_2_15_0[0]), (output_0_3_sva_2_15_0[0]), (output_0_4_sva_2_15_0[0]),
          (output_0_5_sva_2_15_0[0]), (output_0_6_sva_2_15_0[0]), (output_0_7_sva_2_15_0[0]),
          (output_0_8_sva_2_15_0[0]), (output_0_9_sva_2_15_0[0]), (output_0_10_sva_2_15_0[0]),
          (output_0_11_sva_2_15_0[0]), (output_0_12_sva_2_15_0[0]), (output_0_13_sva_2_15_0[0]),
          (output_0_14_sva_2_15_0[0]), (output_0_15_sva_2_15_0[0]), {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
          , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
      strm_out_rsci_idat_31_18 <= MUX_v_14_16_2(output_0_0_sva_2_29_16, output_0_1_sva_2_29_16,
          output_0_2_sva_2_29_16, output_0_3_sva_2_29_16, output_0_4_sva_2_29_16,
          output_0_5_sva_2_29_16, output_0_6_sva_2_29_16, output_0_7_sva_2_29_16,
          output_0_8_sva_2_29_16, output_0_9_sva_2_29_16, output_0_10_sva_2_29_16,
          output_0_11_sva_2_29_16, output_0_12_sva_2_29_16, output_0_13_sva_2_29_16,
          output_0_14_sva_2_29_16, output_0_15_sva_2_29_16, {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
          , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_39 <= 1'b0;
      attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_38_0 <= 39'b000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_3_0_0_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_attn_output_and_4_cse ) begin
      attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2 <= attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2_mx1;
      attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2 <= attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2_mx1;
      attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2 <= attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2_mx1;
      attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2 <= attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2_mx1;
      attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2 <= attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2_mx1;
      attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2 <= attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2_mx1;
      attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2 <= attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2_mx1;
      attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2 <= attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2_mx1;
      attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_39 <= attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_39;
      attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_38_0 <= attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_38_0;
      attention_2_1_16_16_4_4_attn_output_3_0_0_sva_2 <= MUX_v_40_2_2(acc_3_cse_40_1,
          attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3, nand_302_cse);
      attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2 <= attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2_mx1;
      attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2 <= attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2_mx1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_3_0_1_sva_2 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (attention_2_1_16_16_4_4_attn_output_and_13_cse
        | attention_2_1_16_16_4_4_attn_output_and_14_cse) ) begin
      attention_2_1_16_16_4_4_attn_output_3_0_1_sva_2 <= MUX_v_40_2_2(acc_3_cse_40_1,
          attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3, attention_2_1_16_16_4_4_attn_output_and_14_cse);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_3_0_2_sva_2 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (attention_2_1_16_16_4_4_attn_output_and_15_cse
        | attention_2_1_16_16_4_4_attn_output_and_16_cse) ) begin
      attention_2_1_16_16_4_4_attn_output_3_0_2_sva_2 <= MUX_v_40_2_2(acc_3_cse_40_1,
          attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3, attention_2_1_16_16_4_4_attn_output_and_16_cse);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_3_0_3_sva_2 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (attention_2_1_16_16_4_4_attn_output_and_17_cse
        | attention_2_1_16_16_4_4_attn_output_and_18_cse) ) begin
      attention_2_1_16_16_4_4_attn_output_3_0_3_sva_2 <= MUX_v_40_2_2(acc_3_cse_40_1,
          attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3, attention_2_1_16_16_4_4_attn_output_and_18_cse);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_attn_weights_and_36_cse ) begin
      attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2_mx1,
          attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_3, and_dcpl_197);
      attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2_mx1,
          attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_3, and_dcpl_197);
      attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2_mx1,
          attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_3, and_dcpl_197);
      attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2_mx1,
          attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_3, and_dcpl_197);
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2_mx1,
          attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_3, and_dcpl_197);
      attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2_mx1,
          attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_3, and_dcpl_197);
      attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2_mx1,
          attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_3, and_dcpl_197);
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2_mx1,
          attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_3, and_dcpl_197);
      attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2_mx1,
          attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_3, and_dcpl_197);
      attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2_mx1,
          attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_3, and_dcpl_197);
      attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2_mx1,
          attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_3, and_dcpl_197);
      attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2_mx1,
          attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_3, and_dcpl_197);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_2_0_1_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_1_0_1_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_0_0_2_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_2_0_3_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_3_0_0_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_3_0_1_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_3_0_2_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_q_embed_and_5_cse ) begin
      attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1 <= attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1_mx0w1;
      attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1 <= attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1_mx0w1;
      attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1 <= attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1_mx0w1;
      attention_2_1_16_16_4_4_q_embed_2_0_1_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
          attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1, or_dcpl_987);
      attention_2_1_16_16_4_4_q_embed_1_0_1_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
          attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1, or_dcpl_988);
      attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1 <= attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1_mx0w1;
      attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1 <= attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1_mx0w1;
      attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1 <= attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1_mx0w1;
      attention_2_1_16_16_4_4_q_embed_0_0_2_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
          attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1, or_dcpl_996);
      attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1 <= attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1_mx0w1;
      attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1 <= attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1_mx0w1;
      attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1 <= attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1_mx0w1;
      attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1 <= attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1_mx0w1;
      attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1 <= attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1_mx0w1;
      attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1 <= attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1_mx0w1;
      attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1 <= attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1_mx0w1;
      attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1 <= attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1_mx0w1;
      attention_2_1_16_16_4_4_k_embed_2_0_3_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
          attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3, or_dcpl_991);
      attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1 <= attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1_mx0w1;
      attention_2_1_16_16_4_4_k_embed_3_0_0_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
          attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3, or_dcpl_995);
      attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1 <= attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1_mx0w1;
      attention_2_1_16_16_4_4_k_embed_3_0_1_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
          attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3, or_dcpl_997);
      attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1 <= attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1_mx0w1;
      attention_2_1_16_16_4_4_k_embed_3_0_2_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1,
          attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3, or_dcpl_999);
      attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1 <= attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_embed_2_0_3_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_3_0_0_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_3_0_1_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_3_0_2_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_3_0_3_sva_1 <= 40'b0000000000000000000000000000000000000000;
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd <= 1'b0;
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd_1 <= 1'b0;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_47_40
          <= 8'b00000000;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_39
          <= 1'b0;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_38
          <= 1'b0;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_37
          <= 1'b0;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_36
          <= 1'b0;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_35
          <= 1'b0;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_34
          <= 1'b0;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_33
          <= 1'b0;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_32
          <= 1'b0;
      operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_34 <= 1'b0;
      operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_33_0 <= 34'b0000000000000000000000000000000000;
      operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_39 <= 1'b0;
      operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_38_35 <= 4'b0000;
      SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_55 <= 1'b0;
      SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_54_16 <= 39'b000000000000000000000000000000000000000;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_71_48
          <= 24'b000000000000000000000000;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_59_39
          <= 21'b000000000000000000000;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_38_0
          <= 39'b000000000000000000000000000000000000000;
      SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_39 <= 1'b0;
      SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_38_0 <= 39'b000000000000000000000000000000000000000;
      reg_strm_out_rsci_iswt0_cse <= 1'b0;
      reg_strm_in_rsci_iswt0_cse <= 1'b0;
      reg_rms_norm_16_div_cmp_b_ftd_59_38 <= 22'b0000000000000000000000;
      reg_rms_norm_16_div_cmp_b_ftd_37_0 <= 38'b00000000000000000000000000000000000000;
      reg_rms_norm_16_div_cmp_b_ftd_1 <= 1'b0;
      reg_rms_norm_16_div_cmp_a_ftd <= 24'b000000000000000000000000;
      reg_rms_norm_16_div_cmp_a_ftd_1_15_8 <= 8'b00000000;
      reg_rms_norm_16_div_cmp_a_ftd_1_7 <= 1'b0;
      reg_rms_norm_16_div_cmp_a_ftd_1_6 <= 1'b0;
      reg_rms_norm_16_div_cmp_a_ftd_1_5 <= 1'b0;
      reg_rms_norm_16_div_cmp_a_ftd_1_4 <= 1'b0;
      reg_rms_norm_16_div_cmp_a_ftd_1_3 <= 1'b0;
      reg_rms_norm_16_div_cmp_a_ftd_1_2 <= 1'b0;
      reg_rms_norm_16_div_cmp_a_ftd_1_1 <= 1'b0;
      reg_rms_norm_16_div_cmp_a_ftd_1_0 <= 1'b0;
      reg_RMS_NORM_LOOP_1_1_slc_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_mul_55_16_cse_1_slc
          <= 16'b0000000000000000;
      operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_17_16
          <= 2'b00;
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0 <= 1'b0;
      attention_abs_3_qr_sva_38_0 <= 39'b000000000000000000000000000000000000000;
      RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_mux1h_itm <= 1'b0;
      RMS_NORM_LOOP_2_and_29_ssc <= 1'b0;
      RMS_NORM_LOOP_2_and_34_ssc <= 1'b0;
      RMS_NORM_LOOP_2_and_30_m1c <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_8 <= 8'b00000000;
      reg_QUANTIZE_ACTIVATION_LOOP_3_quantized_value_slc_63_32_cse_slc <= 8'b00000000;
      attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0 <= 16'b0000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0 <= 16'b0000000000000000;
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_39_16 <= 24'b000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_39_16 <= 24'b000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_15_8 <= 8'b00000000;
      LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1 <= 1'b0;
      LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_39_16 <= 24'b000000000000000000000000;
      APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm <= 56'b00000000000000000000000000000000000000000000000000000000;
      APPLY_ROTARY_POS_EMB_LOOP_6_mul_3_itm <= 56'b00000000000000000000000000000000000000000000000000000000;
      APPLY_ROTARY_POS_EMB_LOOP_6_mul_itm <= 56'b00000000000000000000000000000000000000000000000000000000;
      APPLY_ROTARY_POS_EMB_LOOP_6_mul_1_itm <= 56'b00000000000000000000000000000000000000000000000000000000;
      TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_16_psp_1 <= 3'b000;
      attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6 <= 40'b0000000000000000000000000000000000000000;
      operator_80_48_true_AC_TRN_AC_WRAP_operator_80_48_true_AC_TRN_AC_WRAP_slc_SOFTMAX_LOOP_4_sqr_56_1_itm_slc
          <= 1'b0;
      attention_abs_5_qr_sva_38_0 <= 39'b000000000000000000000000000000000000000;
      attention_abs_7_qr_sva_38_0 <= 39'b000000000000000000000000000000000000000;
      RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_mux1h_itm <= 1'b0;
      RMS_NORM_LOOP_2_2_and_29_ssc <= 1'b0;
      RMS_NORM_LOOP_2_2_and_34_ssc <= 1'b0;
      RMS_NORM_LOOP_2_2_and_30_m1c <= 1'b0;
      output_0_7_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_7_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_8_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_8_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_6_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_6_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_9_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_9_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_5_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_5_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_10_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_10_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_4_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_4_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_11_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_11_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_3_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_3_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_12_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_12_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_2_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_2_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_13_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_13_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_1_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_1_lpi_3_15_8 <= 8'b00000000;
      output_0_1_lpi_3_7 <= 1'b0;
      output_0_1_lpi_3_6 <= 1'b0;
      output_0_1_lpi_3_5 <= 1'b0;
      output_0_1_lpi_3_4 <= 1'b0;
      output_0_1_lpi_3_3 <= 1'b0;
      output_0_1_lpi_3_2 <= 1'b0;
      output_0_1_lpi_3_1 <= 1'b0;
      output_0_1_lpi_3_0 <= 1'b0;
      output_0_14_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_14_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_0_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_0_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_15_lpi_3_39_16 <= 24'b000000000000000000000000;
      output_0_15_lpi_3_15_0 <= 16'b0000000000000000;
      output_0_15_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_0_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_14_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_1_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_13_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_2_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_12_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_3_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_11_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_4_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_10_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_5_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_9_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_6_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_8_lpi_4_39_16 <= 24'b000000000000000000000000;
      output_0_7_lpi_4_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 ) begin
      attention_2_1_16_16_4_4_q_embed_2_0_3_sva_1 <= attention_2_1_16_16_4_4_q_embed_mux_7_cse;
      attention_2_1_16_16_4_4_q_embed_3_0_0_sva_1 <= attention_2_1_16_16_4_4_q_embed_mux_9_cse;
      attention_2_1_16_16_4_4_q_embed_3_0_1_sva_1 <= attention_2_1_16_16_4_4_q_embed_mux_11_cse;
      attention_2_1_16_16_4_4_q_embed_3_0_2_sva_1 <= attention_2_1_16_16_4_4_q_embed_mux_13_cse;
      attention_2_1_16_16_4_4_q_embed_3_0_3_sva_1 <= attention_2_1_16_16_4_4_q_embed_mux_14_cse;
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd <= mux_816_ssc;
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_a_32_0_ftd_1 <= ~ mux_816_ssc;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_47_40
          <= MUX_v_8_2_2(8'b00000000, operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_nl,
          not_4947_nl);
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_39
          <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_1_nl & (~ or_dcpl_1048);
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_38
          <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_2_nl | or_dcpl_1048;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_37
          <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_3_nl | or_dcpl_1048;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_36
          <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_4_nl | or_dcpl_1048;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_35
          <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_5_nl | or_dcpl_1048;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_34
          <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_6_nl | or_dcpl_1048;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_33
          <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_7_nl | or_dcpl_1048;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_32
          <= operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_8_nl | or_dcpl_1048;
      operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_34 <= MUX1HOT_s_1_7_2(compute_sqrt_guess_sva_34,
          attention_abs_qr_35_0_lpi_1_dfm_mx1_35, (compute_sqrt_for_acc_1_itm_40_1_1[34]),
          (attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_38_0[34]),
          (reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[34]), compute_sqrt_1_guess_sva_34,
          (compute_sqrt_1_for_acc_1_itm_40_1_1[34]), {and_303_ssc , compute_sqrt_guess_or_1_ssc
          , and_dcpl_290 , and_dcpl_276 , and_dcpl_278 , and_315_ssc , and_dcpl_292});
      operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_33_0 <= MUX1HOT_v_34_7_2(compute_sqrt_guess_sva_33_0,
          attention_abs_qr_35_0_lpi_1_dfm_mx1_34_1, (compute_sqrt_for_acc_1_itm_40_1_1[33:0]),
          (attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_38_0[33:0]),
          (reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[33:0]), compute_sqrt_1_guess_sva_33_0,
          (compute_sqrt_1_for_acc_1_itm_40_1_1[33:0]), {and_303_ssc , compute_sqrt_guess_or_1_ssc
          , and_dcpl_290 , and_dcpl_276 , and_dcpl_278 , and_315_ssc , and_dcpl_292});
      operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_39 <= rms_norm_16_mux1h_nl &
          (~ mux_851_ssc);
      operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_b_38_35 <= MUX_v_4_2_2(4'b0000,
          rms_norm_16_mux1h_9_nl, operator_40_24_true_AC_TRN_AC_WRAP_1_not_1_nl);
      SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_55 <= SOFTMAX_LOOP_5_mux_24_nl &
          (~ and_334_ssc);
      SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_a_54_16 <= MUX1HOT_v_39_3_2((SOFTMAX_LOOP_5_mux_12_psp_mx0w0[38:0]),
          reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1, 39'b000000000000000000000010000000000000000,
          {and_dcpl_294 , and_329_ssc , and_334_ssc});
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_a_71_48
          <= MUX_v_24_2_2(24'b000000000000000000000000, LINEAR_FORWARD_NO_MUL_LOOP_2_2_mux1h_2_nl,
          LINEAR_FORWARD_NO_MUL_LOOP_2_2_not_nl);
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_59_39
          <= MUX1HOT_v_21_5_2((z_out_9[59:39]), (LINEAR_FORWARD_NO_MUL_LOOP_2_2_mul_mut[59:39]),
          ({{20{attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_39}},
          attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_39}),
          ({{20{reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd}}, reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd}),
          (LINEAR_FORWARD_NO_MUL_LOOP_2_3_mul_mut[59:39]), {LINEAR_FORWARD_NO_MUL_LOOP_2_2_or_1_cse
          , and_dcpl_260 , and_336_ssc , mux_856_ssc , and_dcpl_268});
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_b_38_0
          <= MUX1HOT_v_39_5_2((z_out_9[38:0]), (LINEAR_FORWARD_NO_MUL_LOOP_2_2_mul_mut[38:0]),
          attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_38_0,
          reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1, (LINEAR_FORWARD_NO_MUL_LOOP_2_3_mul_mut[38:0]),
          {LINEAR_FORWARD_NO_MUL_LOOP_2_2_or_1_cse , and_dcpl_260 , and_336_ssc ,
          mux_856_ssc , and_dcpl_268});
      SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_39 <= MUX1HOT_s_1_3_2((softmax_1_4_3_sum_sva_1[39]),
          (compute_sqrt_1_for_acc_1_itm_40_1_1[39]), reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd,
          {and_dcpl_304 , and_dcpl_292 , and_339_ssc});
      SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_b_38_0 <= MUX1HOT_v_39_3_2((softmax_1_4_3_sum_sva_1[38:0]),
          (compute_sqrt_1_for_acc_1_itm_40_1_1[38:0]), reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1,
          {and_dcpl_304 , and_dcpl_292 , and_339_ssc});
      reg_strm_out_rsci_iswt0_cse <= and_dcpl_306;
      reg_strm_in_rsci_iswt0_cse <= ~(or_1851_cse | (fsm_output[3]) | or_1984_cse
          | mux_862_nl | or_255_cse);
      reg_rms_norm_16_div_cmp_b_ftd_59_38 <= MUX1HOT_v_22_5_2((signext_22_1(compute_sqrt_for_acc_1_itm_40_1_1[39])),
          ({{21{reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd}}, reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd}),
          (LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2[60:39]), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut[60:39]),
          (LINEAR_FORWARD_NO_MUL_LOOP_2_mul_itm[59:38]), {and_dcpl_290 , and_343_itm
          , and_dcpl_257 , and_dcpl_260 , and_dcpl_310});
      reg_rms_norm_16_div_cmp_b_ftd_37_0 <= MUX1HOT_v_38_5_2((compute_sqrt_for_acc_1_itm_40_1_1[38:1]),
          (reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[38:1]), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2[38:1]),
          (LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut[38:1]), (LINEAR_FORWARD_NO_MUL_LOOP_2_mul_itm[37:0]),
          {and_dcpl_290 , and_343_itm , and_dcpl_257 , and_dcpl_260 , and_dcpl_310});
      reg_rms_norm_16_div_cmp_b_ftd_1 <= rms_norm_16_mux1h_10_nl & (~ and_dcpl_310);
      reg_rms_norm_16_div_cmp_a_ftd <= MUX_v_24_2_2(24'b000000000000000000000000,
          rms_norm_16_mux1h_6_nl, rms_norm_16_not_nl);
      reg_rms_norm_16_div_cmp_a_ftd_1_15_8 <= MUX_v_8_2_2(8'b00000000, rms_norm_16_mux1h_7_nl,
          rms_norm_16_not_1_nl);
      reg_rms_norm_16_div_cmp_a_ftd_1_7 <= rms_norm_16_mux1h_11_nl & (~ rms_norm_16_div_cmp_a_mx0c0);
      reg_rms_norm_16_div_cmp_a_ftd_1_6 <= rms_norm_16_mux1h_13_nl & (~ rms_norm_16_div_cmp_a_mx0c0);
      reg_rms_norm_16_div_cmp_a_ftd_1_5 <= rms_norm_16_mux1h_14_nl & (~ rms_norm_16_div_cmp_a_mx0c0);
      reg_rms_norm_16_div_cmp_a_ftd_1_4 <= rms_norm_16_mux1h_15_nl & (~ rms_norm_16_div_cmp_a_mx0c0);
      reg_rms_norm_16_div_cmp_a_ftd_1_3 <= rms_norm_16_mux1h_16_nl & (~ rms_norm_16_div_cmp_a_mx0c0);
      reg_rms_norm_16_div_cmp_a_ftd_1_2 <= rms_norm_16_mux1h_17_nl & (~ rms_norm_16_div_cmp_a_mx0c0);
      reg_rms_norm_16_div_cmp_a_ftd_1_1 <= rms_norm_16_mux1h_18_nl & (~ rms_norm_16_div_cmp_a_mx0c0);
      reg_rms_norm_16_div_cmp_a_ftd_1_0 <= rms_norm_16_mux1h_19_nl | rms_norm_16_div_cmp_a_mx0c0;
      reg_RMS_NORM_LOOP_1_1_slc_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_mul_55_16_cse_1_slc
          <= z_out_10[55:40];
      operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_17_16
          <= operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z[17:16];
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_15_8,
          attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8, and_dcpl_626);
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_7,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_38_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_6,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_39_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_5,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_40_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_4,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_41_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_3,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_42_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_2,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_43_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_1,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_44_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_0,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_15_8,
          attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8, and_dcpl_626);
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_1_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_7,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_24_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_6,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_5,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_26_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_4,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_27_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_3,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_28_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_2,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_29_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_1,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_30_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_0,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_15_8,
          attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8, and_dcpl_626);
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_2_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_7,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_10_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_6,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_11_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_5,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_12_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_4,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_13_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_3,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_14_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_2,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_15_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_1,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_16_nl,
          attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_0,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_15_8,
          attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8, and_dcpl_626);
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_3_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_7,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_17_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_6,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_18_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_5,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_19_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_4,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_20_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_3,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_21_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_2,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_22_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_1,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_23_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_0,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_15_8,
          attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8, and_dcpl_626);
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_4_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_7,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_31_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_6,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_32_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_5,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_33_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_4,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_34_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_3,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_35_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_2,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_36_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_1,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_37_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_0,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_15_8,
          attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8, and_dcpl_626);
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_5_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_7,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_45_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_6,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_46_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_5,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_47_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_4,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_48_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_3,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_49_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_2,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_50_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_1,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_51_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_0,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_15_8,
          attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8, and_dcpl_626);
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_6_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_7,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_52_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_6,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_53_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_5,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_54_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_4,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_55_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_3,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_56_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_2,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_57_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_1,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_58_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_0,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_15_8,
          attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8, and_dcpl_626);
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_7_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_7,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_59_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_6,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_60_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_5,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_61_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_4,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_62_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_3,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_63_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_2,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_64_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_1,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_65_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_0,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_15_8,
          attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8, and_dcpl_626);
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_8_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_7,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_66_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_6,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_67_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_5,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_68_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_4,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_69_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_3,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_70_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_2,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_71_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_1,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_72_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_0,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_15_8,
          attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8, and_dcpl_626);
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_9_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_7,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_73_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_6,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_74_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_5,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_75_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_4,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_76_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_3,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_77_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_2,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_78_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_1,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0 <= MUX1HOT_s_1_3_2(INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_79_nl,
          attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_0,
          {and_dcpl_622 , and_dcpl_240 , and_dcpl_626});
      attention_abs_3_qr_sva_38_0 <= attention_abs_2_mux_2[38:0];
      RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_mux1h_itm <= MUX1HOT_s_1_3_2((attention_abs_1_qr_sva_1[39]),
          reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1, (attention_abs_2_mux_2[39]),
          {and_28_cse , RMS_NORM_LOOP_2_and_29_ssc_1 , RMS_NORM_LOOP_2_and_34_ssc_1});
      RMS_NORM_LOOP_2_and_29_ssc <= RMS_NORM_LOOP_2_and_29_ssc_1;
      RMS_NORM_LOOP_2_and_34_ssc <= RMS_NORM_LOOP_2_and_34_ssc_1;
      RMS_NORM_LOOP_2_and_30_m1c <= RMS_NORM_LOOP_2_and_30_m1c_1;
      attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_15_8,
          attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8, and_dcpl_626);
      reg_QUANTIZE_ACTIVATION_LOOP_3_quantized_value_slc_63_32_cse_slc <= z_out_10[63:56];
      attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_5_nl, not_4472_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_30_nl, not_4469_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_32_nl, not_4468_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_34_nl, not_4467_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_36_nl, not_4466_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_38_nl, not_4465_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_42_nl, not_4463_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_44_nl, not_4462_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_46_nl, not_4461_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_48_nl, not_4460_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_50_nl, not_4459_nl);
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          ({attention_2_1_16_16_4_4_k_proj_re_mux1h_68_nl , attention_2_1_16_16_4_4_k_proj_re_mux1h_118_nl}),
          not_4443_nl);
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_58_nl, not_4582_nl);
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_59_nl, not_4583_nl);
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_60_nl, not_4584_nl);
      attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_61_nl, not_4585_nl);
      attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_62_nl, not_4586_nl);
      attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_63_nl, not_4587_nl);
      attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_64_nl, not_4588_nl);
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_15_8 <= MUX_v_8_2_2(attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_15_8,
          attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8, and_dcpl_626);
      LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_1 <= (LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_2[1])
          & (~ mux_2100_ssc);
      LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0 <= QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_1_nl
          & (~ mux_2100_ssc);
      attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16 <= MUX_v_24_2_2(apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_39_16,
          attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16 <= MUX_v_24_2_2(LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48,
          attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16 <= MUX_v_24_2_2(apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_39_16,
          attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16 <= MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_39_16,
          attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16 <= MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16,
          attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_39_16,
          attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16 <= MUX_v_24_2_2(for_for_strm_in_tmp_sva_25_2,
          attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16,
          attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_39_16,
          attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_39_16,
          attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_39_16,
          attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16 <= MUX_v_24_2_2(apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16 <= MUX_v_24_2_2(apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_3_39_16,
          attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16 <= MUX_v_24_2_2(apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16 <= MUX_v_24_2_2(apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16 <= MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_3_39_16,
          attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16_mx1, and_dcpl_725);
      attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_39_16 <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16,
          attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16_mx0w1,
          attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16, {and_dcpl_1073 , and_dcpl_240
          , and_dcpl_207 , and_dcpl_847});
      attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_39_16 <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16,
          attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16_mx0w1,
          attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16, {and_dcpl_1073 , and_dcpl_240
          , and_dcpl_207 , and_dcpl_847});
      attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_39_16 <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16,
          attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16_mx0w1,
          attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16, {and_dcpl_1073 , and_dcpl_240
          , and_dcpl_207 , and_dcpl_847});
      attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_39_16 <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16,
          attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16,
          attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16_mx0w1, {operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse
          , and_dcpl_240 , attention_2_1_16_16_4_4_k_proj_re_or_17_cse , and_dcpl_207});
      attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_39_16 <= MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16,
          attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16_mx0w1,
          attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16, {and_dcpl_1073 , and_dcpl_240
          , and_dcpl_207 , and_dcpl_847});
      APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm <= z_out_10[55:0];
      APPLY_ROTARY_POS_EMB_LOOP_6_mul_3_itm <= nl_APPLY_ROTARY_POS_EMB_LOOP_6_mul_3_itm[55:0];
      APPLY_ROTARY_POS_EMB_LOOP_6_mul_itm <= $unsigned(nl_APPLY_ROTARY_POS_EMB_LOOP_6_mul_sgnd);
      APPLY_ROTARY_POS_EMB_LOOP_6_mul_1_itm <= z_out_9[55:0];
      TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_16_psp_1 <= nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_16_psp_1[2:0];
      attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2,
          attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_3,
          {and_dcpl_1193 , and_dcpl_1194 , and_dcpl_1195});
      attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2,
          attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_3,
          {and_dcpl_1193 , and_dcpl_1194 , and_dcpl_1195});
      attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2,
          attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_3,
          {and_dcpl_1193 , and_dcpl_1194 , and_dcpl_1195});
      attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2,
          attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_3,
          {and_dcpl_1193 , and_dcpl_1194 , and_dcpl_1195});
      attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2,
          attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_3,
          {and_dcpl_1193 , and_dcpl_1194 , and_dcpl_1195});
      attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2,
          attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_3,
          {and_dcpl_1193 , and_dcpl_1194 , and_dcpl_1195});
      attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2,
          attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_3,
          {and_dcpl_1193 , and_dcpl_1194 , and_dcpl_1195});
      attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2,
          attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_3,
          {and_dcpl_1193 , and_dcpl_1194 , and_dcpl_1195});
      attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2,
          attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_3,
          {and_dcpl_1193 , and_dcpl_1194 , and_dcpl_1195});
      attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2,
          attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_3,
          {and_dcpl_1193 , and_dcpl_1194 , and_dcpl_1195});
      attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2,
          attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_3,
          {and_dcpl_1193 , and_dcpl_1194 , and_dcpl_1195});
      attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6 <= MUX1HOT_v_40_3_2(attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2,
          attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6_mx1, attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_3,
          {and_dcpl_1193 , and_dcpl_1194 , and_dcpl_1195});
      operator_80_48_true_AC_TRN_AC_WRAP_operator_80_48_true_AC_TRN_AC_WRAP_slc_SOFTMAX_LOOP_4_sqr_56_1_itm_slc
          <= z_out_10[56];
      attention_abs_5_qr_sva_38_0 <= attention_abs_5_qr_sva_1[38:0];
      attention_abs_7_qr_sva_38_0 <= attention_abs_6_mux_2[38:0];
      RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_mux1h_itm <= MUX1HOT_s_1_3_2((attention_abs_5_qr_sva_1[39]),
          reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1, (attention_abs_6_mux_2[39]),
          {RMS_NORM_LOOP_2_2_and_32_ssc_mx0w3 , RMS_NORM_LOOP_2_2_and_29_ssc_1 ,
          RMS_NORM_LOOP_2_2_and_34_ssc_1});
      RMS_NORM_LOOP_2_2_and_29_ssc <= RMS_NORM_LOOP_2_2_and_29_ssc_1;
      RMS_NORM_LOOP_2_2_and_34_ssc <= RMS_NORM_LOOP_2_2_and_34_ssc_1;
      RMS_NORM_LOOP_2_2_and_30_m1c <= RMS_NORM_LOOP_2_2_and_30_m1c_1;
      output_0_7_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_nl,
          not_4589_nl);
      output_0_7_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_44_nl,
          not_4590_nl);
      output_0_8_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_36_nl,
          not_4591_nl);
      output_0_8_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_45_nl,
          not_4592_nl);
      output_0_6_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_37_nl,
          not_4593_nl);
      output_0_6_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_46_nl,
          not_4594_nl);
      output_0_9_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_38_nl,
          not_4595_nl);
      output_0_9_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_47_nl,
          not_4596_nl);
      output_0_5_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_39_nl,
          not_4597_nl);
      output_0_5_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_48_nl,
          not_4598_nl);
      output_0_10_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_40_nl,
          not_4599_nl);
      output_0_10_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_49_nl,
          not_4600_nl);
      output_0_4_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_41_nl,
          not_4601_nl);
      output_0_4_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_50_nl,
          not_4602_nl);
      output_0_11_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_42_nl,
          not_4603_nl);
      output_0_11_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_51_nl,
          not_4604_nl);
      output_0_3_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_43_nl,
          not_4605_nl);
      output_0_3_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_52_nl,
          not_4606_nl);
      output_0_12_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_44_nl,
          not_4607_nl);
      output_0_12_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_53_nl,
          not_4608_nl);
      output_0_2_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_45_nl,
          not_4609_nl);
      output_0_2_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_54_nl,
          not_4610_nl);
      output_0_13_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_46_nl,
          not_4611_nl);
      output_0_13_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_55_nl,
          not_4612_nl);
      output_0_1_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_47_nl,
          not_4613_nl);
      output_0_1_lpi_3_15_8 <= MUX_v_8_2_2(8'b00000000, attention_2_1_16_16_4_4_k_proj_re_mux_56_nl,
          not_5055_nl);
      output_0_1_lpi_3_7 <= attention_2_1_16_16_4_4_k_proj_re_mux_60_nl & (~ and_dcpl_1154);
      output_0_1_lpi_3_6 <= attention_2_1_16_16_4_4_k_proj_re_mux_61_nl & (~ and_dcpl_1154);
      output_0_1_lpi_3_5 <= attention_2_1_16_16_4_4_k_proj_re_mux_62_nl & (~ and_dcpl_1154);
      output_0_1_lpi_3_4 <= attention_2_1_16_16_4_4_k_proj_re_mux_63_nl & (~ and_dcpl_1154);
      output_0_1_lpi_3_3 <= attention_2_1_16_16_4_4_k_proj_re_mux_64_nl & (~ and_dcpl_1154);
      output_0_1_lpi_3_2 <= attention_2_1_16_16_4_4_k_proj_re_mux_65_nl & (~ and_dcpl_1154);
      output_0_1_lpi_3_1 <= attention_2_1_16_16_4_4_k_proj_re_mux_66_nl & (~ and_dcpl_1154);
      output_0_1_lpi_3_0 <= attention_2_1_16_16_4_4_k_proj_re_mux_67_nl & (~ and_dcpl_1154);
      output_0_14_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_48_nl,
          not_4615_nl);
      output_0_14_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_57_nl,
          not_4616_nl);
      output_0_0_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_49_nl,
          not_4617_nl);
      output_0_0_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_58_nl,
          not_4618_nl);
      output_0_15_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000, attention_2_1_16_16_4_4_v_proj_re_mux_50_nl,
          not_4619_nl);
      output_0_15_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000, attention_2_1_16_16_4_4_k_proj_re_mux_59_nl,
          not_4620_nl);
      output_0_15_lpi_4_39_16 <= MUX_v_24_2_2(output_0_15_lpi_3_39_16, output_0_15_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_0_lpi_4_39_16 <= MUX_v_24_2_2(output_0_0_lpi_3_39_16, output_0_0_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_14_lpi_4_39_16 <= MUX_v_24_2_2(output_0_14_lpi_3_39_16, output_0_14_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_1_lpi_4_39_16 <= MUX_v_24_2_2(output_0_1_lpi_3_39_16, output_0_1_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_13_lpi_4_39_16 <= MUX_v_24_2_2(output_0_13_lpi_3_39_16, output_0_13_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_2_lpi_4_39_16 <= MUX_v_24_2_2(output_0_2_lpi_3_39_16, output_0_2_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_12_lpi_4_39_16 <= MUX_v_24_2_2(output_0_12_lpi_3_39_16, output_0_12_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_3_lpi_4_39_16 <= MUX_v_24_2_2(output_0_3_lpi_3_39_16, output_0_3_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_11_lpi_4_39_16 <= MUX_v_24_2_2(output_0_11_lpi_3_39_16, output_0_11_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_4_lpi_4_39_16 <= MUX_v_24_2_2(output_0_4_lpi_3_39_16, output_0_4_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_10_lpi_4_39_16 <= MUX_v_24_2_2(output_0_10_lpi_3_39_16, output_0_10_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_5_lpi_4_39_16 <= MUX_v_24_2_2(output_0_5_lpi_3_39_16, output_0_5_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_9_lpi_4_39_16 <= MUX_v_24_2_2(output_0_9_lpi_3_39_16, output_0_9_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_6_lpi_4_39_16 <= MUX_v_24_2_2(output_0_6_lpi_3_39_16, output_0_6_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_8_lpi_4_39_16 <= MUX_v_24_2_2(output_0_8_lpi_3_39_16, output_0_8_lpi_4_39_16_mx1,
          and_dcpl_1227);
      output_0_7_lpi_4_39_16 <= MUX_v_24_2_2(output_0_7_lpi_3_39_16, output_0_7_lpi_4_39_16_mx1,
          and_dcpl_1227);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0 <= 16'b0000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16 <= 24'b000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_8 <= 8'b00000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_7 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_6 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_5 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_4 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_3 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_2 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_1 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_0 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16 <= 24'b000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_13 <= 3'b000;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_12_8 <= 5'b00000;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_7 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_6 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_5 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_4 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_3 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_2 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_1 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_0 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16 <= 24'b000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_8 <= 8'b00000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_7 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_6 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_5 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_4 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_3 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_2 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_1 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_0 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_39_16 <= 24'b000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_8 <= 8'b00000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_7 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_6 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_5 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_4 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_3 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_2 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_1 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_0 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16 <= 24'b000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_8 <= 8'b00000000;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_1 <=
          1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_2 <=
          1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_3 <=
          1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_4 <=
          1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_5 <=
          1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_6 <=
          1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_7 <=
          1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16 <= 24'b000000000000000000000000;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_ftd <= 8'b00000000;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_1 <=
          1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_2 <=
          1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_3 <=
          1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_4 <=
          1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_5 <=
          1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_6 <=
          1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_7 <=
          1'b0;
    end
    else if ( attention_2_1_16_16_4_4_v_proj_and_2_cse ) begin
      attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_15_0 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
          attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0, or_dcpl_1010);
      attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_15_0 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
          attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0, or_dcpl_1012);
      attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_15_0 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
          attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0, or_dcpl_1014);
      attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_15_0 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
          attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0, or_dcpl_1016);
      attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_15_0 <= MUX_v_16_2_2(RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
          attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0, or_dcpl_1018);
      attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0 <= attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0_mx0w1;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16_mx0w1;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_8 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_7 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_6 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_5 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_4 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_3 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_2 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_1 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_0 <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16_mx0w1;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_13 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_13;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_12_8 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_12_8;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_7 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_6 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_5 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_4 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_3 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_2 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_1 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_0 <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16_mx0w1;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_8 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_7 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_6 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_5 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_4 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_3 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_2 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_1 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_0 <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_39_16 <= MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1,
          for_for_strm_in_tmp_sva_25_2, or_dcpl_1023);
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_8 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_7 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_6 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_5 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_4 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_3 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_2 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_1 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_0 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16 <= apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16_mx0w1;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_8 <= apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd <= apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_1 <=
          apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_2 <=
          apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_3 <=
          apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_4 <=
          apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_5 <=
          apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_6 <=
          apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_7 <=
          apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16 <= apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16_mx0w1;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_ftd <= apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd <= apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_1 <=
          apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_2 <=
          apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_3 <=
          apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_4 <=
          apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_5 <=
          apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_6 <=
          apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1;
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_7 <=
          apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2 <= 40'b0000000000000000000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2 <= 40'b0000000000000000000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2 <= 40'b0000000000000000000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2 <= 40'b0000000000000000000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( apply_rotary_pos_emb_1_4_4_rotated_q_and_cse ) begin
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2 <= MUX1HOT_v_40_7_2(apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm,
          apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2_mx0w1, attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1,
          attention_2_1_16_16_4_4_k_embed_1_0_0_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2,
          GEMM_3D_FLOAT_LOOP_3_1_and_32_nl, attention_2_1_16_16_4_4_attn_output_1_0_1_sva_2_mx1,
          {apply_rotary_pos_emb_1_4_4_rotated_q_or_11_cse , and_dcpl_207 , apply_rotary_pos_emb_1_4_4_rotated_q_or_12_cse
          , and_dcpl_204 , and_dcpl_220 , and_dcpl_222 , and_dcpl_187});
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2 <= MUX1HOT_v_40_7_2(apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm,
          apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2_mx0w1, attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1,
          attention_2_1_16_16_4_4_k_embed_0_0_3_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2,
          GEMM_3D_FLOAT_LOOP_3_1_and_34_nl, attention_2_1_16_16_4_4_attn_output_1_0_0_sva_2_mx1,
          {apply_rotary_pos_emb_1_4_4_rotated_q_or_11_cse , and_dcpl_207 , apply_rotary_pos_emb_1_4_4_rotated_q_or_12_cse
          , and_dcpl_204 , and_dcpl_220 , and_dcpl_222 , and_dcpl_187});
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2 <= MUX1HOT_v_40_7_2(apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm,
          apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2_mx0w1, attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1,
          attention_2_1_16_16_4_4_k_embed_1_0_1_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2,
          GEMM_3D_FLOAT_LOOP_3_1_and_30_nl, attention_2_1_16_16_4_4_attn_output_1_0_2_sva_2_mx1,
          {apply_rotary_pos_emb_1_4_4_rotated_q_or_11_cse , and_dcpl_207 , apply_rotary_pos_emb_1_4_4_rotated_q_or_12_cse
          , and_dcpl_204 , and_dcpl_220 , and_dcpl_222 , and_dcpl_187});
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2 <= MUX1HOT_v_40_7_2(apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm,
          apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2_mx0w1, attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1,
          attention_2_1_16_16_4_4_k_embed_0_0_1_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2,
          GEMM_3D_FLOAT_LOOP_3_1_and_40_nl, attention_2_1_16_16_4_4_attn_output_0_0_1_sva_2_mx1,
          {apply_rotary_pos_emb_1_4_4_rotated_q_or_11_cse , and_dcpl_207 , apply_rotary_pos_emb_1_4_4_rotated_q_or_12_cse
          , and_dcpl_204 , and_dcpl_220 , and_dcpl_222 , and_dcpl_187});
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2 <= MUX1HOT_v_40_7_2(apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm,
          apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2_mx0w1, attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1,
          attention_2_1_16_16_4_4_k_embed_0_0_2_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2,
          GEMM_3D_FLOAT_LOOP_3_1_and_38_nl, attention_2_1_16_16_4_4_attn_output_0_0_2_sva_2_mx1,
          {apply_rotary_pos_emb_1_4_4_rotated_q_or_11_cse , and_dcpl_207 , apply_rotary_pos_emb_1_4_4_rotated_q_or_12_cse
          , and_dcpl_204 , and_dcpl_220 , and_dcpl_222 , and_dcpl_187});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~(mux_797_nl &
        (~ (fsm_output[8])))) ) begin
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2 <= MUX1HOT_v_40_6_2(apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w0,
          apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w3,
          attention_2_1_16_16_4_4_k_embed_0_0_0_sva_1, GEMM_3D_FLOAT_LOOP_3_1_and_42_nl,
          acc_3_cse_40_1, {and_dcpl_207 , and_259_nl , and_dcpl_204 , and_dcpl_216
          , and_dcpl_222 , and_267_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1028)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_15 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_14_12 <= 3'b000;
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_11_9 <= 3'b000;
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_8 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_13 <= 3'b000;
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0 <= 13'b0000000000000;
      attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_ftd <= 8'b00000000;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd <= 1'b0;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_1 <= 1'b0;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_2 <= 1'b0;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_3 <= 1'b0;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_4 <= 1'b0;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_5 <= 1'b0;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_6 <= 1'b0;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_7 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_8 <= 8'b00000000;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd <= 1'b0;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_1 <= 1'b0;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_2 <= 1'b0;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_3 <= 1'b0;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_4 <= 1'b0;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_5 <= 1'b0;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_6 <= 1'b0;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_7 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_7 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_6 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_5 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_4 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_3 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_2 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_1 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_0 <= 1'b0;
      attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_q_proj_and_23_cse ) begin
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_15_8;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_7;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_6;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_5;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_4;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_3;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_2;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_1;
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_15_8;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_7;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_6;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_5;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_4;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_3;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_2;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_1;
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_15_8;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_7;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_6;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_5;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_4;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_3;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_2;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_1;
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_15_8;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_7;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_6;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_5;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_4;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_3;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_2;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_1;
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_15_8;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_7;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_6;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_5;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_4;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_3;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_2;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_1;
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_15_8;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_7;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_6;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_5;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_4;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_3;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_2;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_1;
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_15_8;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_7;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_6;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_5;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_4;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_3;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_2;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_1;
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_15_8;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_7;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_6;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_5;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_4;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_3;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_2;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_1;
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_15 <= MUX_s_1_2_2((z_out[15]), operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_15,
          or_dcpl_1040);
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_14_12 <= MUX_v_3_2_2((z_out[14:12]),
          reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd,
          or_dcpl_1040);
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_11_9 <= MUX_v_3_2_2((z_out[11:9]),
          reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1,
          or_dcpl_1040);
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_8 <= MUX_s_1_2_2((z_out[8]), reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2,
          or_dcpl_1040);
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0 <= MUX_v_8_2_2((z_out[7:0]),
          reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3,
          or_dcpl_1040);
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_15_8;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_7;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_6;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_5;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_4;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_3;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_2;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_1;
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0 <= attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_15_8;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_7;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_6;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_5;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_4;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_3;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_2;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_1;
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0 <= attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_15_8;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_7;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_6;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_5;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_4;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_3;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_2;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_1;
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_15_8;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_7 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_7;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_6 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_6;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_5 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_5;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_4 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_4;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_3 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_3;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_2 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_2;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_1 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_1;
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_0 <= attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_8 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_15_8;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_7 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_7;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_6 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_6;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_5 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_5;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_4 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_4;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_3 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_3;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_2 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_2;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_1 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_1;
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_0 <= attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_13 <= attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_15_13;
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0 <= attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0;
      attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_15_8 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_13_cse;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_7 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_7;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_6 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_6;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_5 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_5;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_4 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_4;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_3 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_3;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_2 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_2;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_1 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_1;
      attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_0 <= RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_0;
      attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16_mx0w1;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_ftd <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_15_8;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_7;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_1 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_6;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_2 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_5;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_3 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_4;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_4 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_3;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_5 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_2;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_6 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_1;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_7 <= attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_8 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_15_8;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_7;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_1 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_6;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_2 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_5;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_3 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_4;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_4 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_3;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_5 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_2;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_6 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_1;
      reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_7 <= attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_39_16 <= MUX_v_24_2_2(RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
          for_for_strm_in_tmp_sva_25_2, or_dcpl_1017);
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_8 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_15_8;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_7 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_7;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_6 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_6;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_5 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_5;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_4 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_4;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_3 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_3;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_2 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_2;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_1 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_1;
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_0 <= attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_0;
      attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0_mx0w1;
      attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16_mx0w1;
      attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1030)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1031)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1033)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1035)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1037)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1038)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1039)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1040)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1041)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1042)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1043)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1044)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1045)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ or_dcpl_1046)
        & and_dcpl_240 ) begin
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_0_14_sva_1 <= 40'b0000000000000000000000000000000000000000;
      input_0_1_sva_1 <= 40'b0000000000000000000000000000000000000000;
      input_0_13_sva_1_39 <= 1'b0;
      input_0_13_sva_1_38_0 <= 39'b000000000000000000000000000000000000000;
      input_0_2_sva_1_39 <= 1'b0;
      input_0_2_sva_1_38_0 <= 39'b000000000000000000000000000000000000000;
      input_0_12_sva_1 <= 40'b0000000000000000000000000000000000000000;
      input_0_3_sva_1 <= 40'b0000000000000000000000000000000000000000;
      input_0_11_sva_1 <= 40'b0000000000000000000000000000000000000000;
      input_0_4_sva_1 <= 40'b0000000000000000000000000000000000000000;
      input_0_10_sva_1 <= 40'b0000000000000000000000000000000000000000;
      input_0_5_sva_1 <= 40'b0000000000000000000000000000000000000000;
      input_0_9_sva_1 <= 40'b0000000000000000000000000000000000000000;
      input_0_6_sva_1 <= 40'b0000000000000000000000000000000000000000;
      input_0_8_sva_1 <= 40'b0000000000000000000000000000000000000000;
      input_0_7_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( input_and_cse ) begin
      input_0_14_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3,
          input_0_14_sva_2, and_dcpl_248);
      input_0_1_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3,
          input_0_1_sva_2, and_dcpl_248);
      input_0_13_sva_1_39 <= MUX_s_1_2_2(reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd,
          input_0_13_sva_2_39, and_dcpl_248);
      input_0_13_sva_1_38_0 <= MUX_v_39_2_2(reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1,
          input_0_13_sva_2_38_0, and_dcpl_248);
      input_0_2_sva_1_39 <= MUX_s_1_2_2(QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39,
          input_0_2_sva_2_39, and_dcpl_248);
      input_0_2_sva_1_38_0 <= MUX_v_39_2_2(QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0,
          input_0_2_sva_2_38_0, and_dcpl_248);
      input_0_12_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1,
          input_0_12_sva_2, and_dcpl_248);
      input_0_3_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3,
          input_0_3_sva_2, and_dcpl_248);
      input_0_11_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3,
          input_0_11_sva_2, and_dcpl_248);
      input_0_4_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3,
          input_0_4_sva_2, and_dcpl_248);
      input_0_10_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3,
          input_0_10_sva_2, and_dcpl_248);
      input_0_5_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3,
          input_0_5_sva_2, and_dcpl_248);
      input_0_9_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3,
          input_0_9_sva_2, and_dcpl_248);
      input_0_6_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3,
          input_0_6_sva_2, and_dcpl_248);
      input_0_8_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm, input_0_8_sva_2,
          and_dcpl_248);
      input_0_7_sva_1 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1,
          input_0_7_sva_2, and_dcpl_248);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm <= 40'b0000000000000000000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm <= 40'b0000000000000000000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm <= 40'b0000000000000000000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm <= 40'b0000000000000000000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm <= 40'b0000000000000000000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( apply_rotary_pos_emb_1_4_4_rotated_q_and_3_cse ) begin
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm <= apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2_mx0w1;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm <= apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2_mx0w1;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm <= apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2_mx0w1;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm <= apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2_mx0w1;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w0;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm <= apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_15_8 <= 8'b00000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_7 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_6 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_5 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_4 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_3 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_2 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_1 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_0 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd <= 8'b00000000;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_1 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_2 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_3 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_4 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_5 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_6 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_7 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_8 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_39_16 <= 24'b000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_39_16 <= 24'b000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3 <= 40'b0000000000000000000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( apply_rotary_pos_emb_1_4_4_rotated_k_and_6_cse ) begin
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_15_8 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_7 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_6 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_5 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_4 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_2 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_1 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_0 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_1 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_2 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_4 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_5 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_6 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_7 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_8 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_39_16 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_39_16 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1;
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1;
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_15_8 <= 8'b00000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_7 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_6 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_5 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_4 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_3 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_2 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_1 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_0 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd <= 8'b00000000;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_1 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_2 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_3 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_4 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_5 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_6 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_7 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_8 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_39_16 <= 24'b000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_39_16 <= 24'b000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3 <= 40'b0000000000000000000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( apply_rotary_pos_emb_1_4_4_rotated_k_and_7_cse ) begin
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_15_8 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_7 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_6 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_5 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_4 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_2 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_1 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_0 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_1 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_2 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_4 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_5 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_6 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_7 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_8 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_39_16 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_39_16 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1;
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1;
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_15_8 <= 8'b00000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_7 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_6 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_5 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_4 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_3 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_2 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_1 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_0 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd <= 8'b00000000;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_1 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_2 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_3 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_4 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_5 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_6 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_7 <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_8 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_39_16 <= 24'b000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_39_16 <= 24'b000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3 <= 40'b0000000000000000000000000000000000000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( apply_rotary_pos_emb_1_4_4_rotated_k_and_8_cse ) begin
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_15_8 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_7 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_6 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_5 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_4 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_2 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_1 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_0 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_1 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_2 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_4 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_5 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_6 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_7 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_8 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_39_16 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_39_16 <= APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1;
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3 <= APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (((~ or_dcpl_1025)
        & mux_902_nl) | attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c0 |
        and_dcpl_344 | and_dcpl_346 | and_dcpl_204 | and_dcpl_348 | and_dcpl_349
        | and_dcpl_351 | attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c9)
        ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1 <= MUX1HOT_v_40_9_2(({{10{strm_in_rsci_idat_mxwt[29]}},
          strm_in_rsci_idat_mxwt}), input_0_0_sva_2, attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1,
          attention_2_1_16_16_4_4_k_embed_3_0_3_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2,
          attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx1, attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx2,
          ({ATTN_2D_LOOP_3_mux_16_itm , ATTN_2D_LOOP_3_mux_17_itm}), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
          {attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c0 , and_dcpl_344
          , and_dcpl_346 , and_dcpl_204 , and_dcpl_348 , and_dcpl_349 , and_dcpl_351
          , and_dcpl_352 , attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx0c9});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd <= 1'b0;
      reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1 <= 39'b000000000000000000000000000000000000000;
    end
    else if ( GEMM_3D_FLOAT_LOOP_4_1_and_ssc ) begin
      reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd <= rms_norm_16_variance_mux1h_nl & GEMM_3D_FLOAT_LOOP_4_1_nand_itm;
      reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1 <= MUX_v_39_2_2(39'b000000000000000000000000000000000000000,
          rms_norm_16_variance_mux1h_1_nl, GEMM_3D_FLOAT_LOOP_4_1_nand_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd <= 1'b0;
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 <= 1'b0;
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2 <= 2'b00;
    end
    else if ( LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_ssc ) begin
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd <= LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux_nl
          & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_5_itm;
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 <= LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_8_nl
          & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_5_itm;
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2 <= MUX_v_2_2_2(2'b00,
          LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_9_nl, LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_5_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd <= 1'b0;
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 <= 2'b00;
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 <= 1'b0;
    end
    else if ( LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_and_ssc ) begin
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd <= ~((~(compute_sqrt_for_i_mux1h_nl
          & (~ LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c3))) | LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c0);
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 <= ~(MUX_v_2_2_2(compute_sqrt_for_i_nand_1_nl,
          2'b11, LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c0));
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 <= ~((~(compute_sqrt_for_i_mux1h_2_nl
          | LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c3)) | LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c0);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_strm_in_tmp_sva_31_26 <= 6'b000000;
      for_for_strm_in_tmp_sva_25_2 <= 24'b000000000000000000000000;
    end
    else if ( for_for_and_13_ssc ) begin
      for_for_strm_in_tmp_sva_31_26 <= strm_in_rsci_idat_mxwt[29:24];
      for_for_strm_in_tmp_sva_25_2 <= MUX_v_24_2_2((strm_in_rsci_idat_mxwt[23:0]),
          INIT_2D_MEM_LOOP_2_1_and_nl, for_for_strm_in_tmp_sva_31_2_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_1068)
        | GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c0 | GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c1
        | GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c2 | GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c4
        | and_dcpl_313 | GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c7 | and_dcpl_316 |
        GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c9 | GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c10)
        & (mux_1063_nl | (fsm_output[8])) ) begin
      GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm <= MUX1HOT_v_40_10_2(({{10{strm_in_rsci_idat_mxwt[29]}},
          strm_in_rsci_idat_mxwt}), input_0_8_sva_1, rms_norm_16_div_cmp_z_oreg,
          operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z, APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1,
          GEMM_3D_FLOAT_LOOP_4_mux_17_nl, SOFTMAX_LOOP_4_x_acc_2_nl, GEMM_3D_FLOAT_LOOP_4_1_mux_18_nl,
          z_out_2, (SOFTMAX_LOOP_5_SOFTMAX_LOOP_5_div_1_cmp_z[39:0]), {GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c0
          , GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c1 , GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c2
          , GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c4 , and_dcpl_207 , and_dcpl_313
          , GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c7 , and_dcpl_316 , GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c9
          , GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm_mx0c10});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39 <= 1'b0;
      QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0 <= 39'b000000000000000000000000000000000000000;
    end
    else if ( QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_and_ssc ) begin
      QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39 <= MUX1HOT_s_1_13_2((strm_in_rsci_idat_mxwt[29]),
          input_0_2_sva_1_39, RMS_NORM_LOOP_2_mux_22_nl, QUANTIZE_ACTIVATION_LOOP_3_quantized_value_mux_nl,
          (APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1[39]), (attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d[39]),
          (attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1[39]), (attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1[39]),
          (attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1[39]), (attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1[39]),
          (SOFTMAX_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_cse_sva_1[39]),
          (attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d[39]), (z_out_2[39]), {and_474_rgt
          , and_476_rgt , and_dcpl_438 , and_dcpl_439 , and_dcpl_374 , and_480_rgt
          , for_for_and_14_rgt , for_for_and_15_rgt , for_for_and_16_rgt , for_for_and_17_rgt
          , and_485_rgt , and_486_rgt , for_for_or_1_rgt});
      QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0 <= MUX1HOT_v_39_13_2(({{9{strm_in_rsci_idat_mxwt[29]}},
          strm_in_rsci_idat_mxwt}), input_0_2_sva_1_38_0, RMS_NORM_LOOP_2_mux_24_nl,
          QUANTIZE_ACTIVATION_LOOP_3_quantized_value_mux_1_nl, (APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1[38:0]),
          (attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d[38:0]), (attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1[38:0]),
          (attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1[38:0]), (attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1[38:0]),
          (attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1[38:0]), (SOFTMAX_LOOP_3_slc_attention_2_1_16_16_4_4_attn_weights_40_39_0_cse_sva_1[38:0]),
          (attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d[38:0]), (z_out_2[38:0]),
          {and_474_rgt , and_476_rgt , and_dcpl_438 , and_dcpl_439 , and_dcpl_374
          , and_480_rgt , for_for_and_14_rgt , for_for_and_15_rgt , for_for_and_16_rgt
          , for_for_and_17_rgt , and_485_rgt , and_486_rgt , for_for_or_1_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_998)
        | attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c0 | attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c1
        | (~ mux_1079_itm) | and_dcpl_204 | and_dcpl_216 | and_dcpl_348 | and_dcpl_351
        | attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c7 | attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c9)
        ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          for_for_mux1h_5_nl, attention_2_1_16_16_4_4_attn_output_2D_not_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_989)
        | attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c0 | attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c1
        | and_dcpl_346 | (~ mux_1099_nl) | and_dcpl_204 | and_dcpl_348 | and_dcpl_351
        | attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c7 | attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c9)
        & (attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c0 | attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c1
        | and_dcpl_346 | and_dcpl_204 | and_dcpl_348 | and_dcpl_351 | attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c7
        | and_dcpl_352 | attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c9)
        ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          for_for_mux1h_6_nl, attention_2_1_16_16_4_4_attn_output_2D_not_3_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd <= 1'b0;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1 <= 39'b000000000000000000000000000000000000000;
    end
    else if ( apply_rotary_pos_emb_1_4_4_rotated_q_and_37_cse ) begin
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd <= MUX1HOT_s_1_6_2((strm_in_rsci_idat_mxwt[29]),
          input_0_13_sva_1_39, (APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1[39]),
          attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_39, GEMM_3D_FLOAT_LOOP_3_1_and_36_nl,
          attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_39, {apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c0
          , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c1 , and_dcpl_207
          , and_dcpl_220 , and_dcpl_222 , and_dcpl_187});
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1 <= MUX1HOT_v_39_8_2(({{9{strm_in_rsci_idat_mxwt[29]}},
          strm_in_rsci_idat_mxwt}), input_0_13_sva_1_38_0, QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_dfm_1_38_0_1,
          QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_dfm_1_38_0_mx0w1, (APPLY_ROTARY_POS_EMB_LOOP_3_acc_6_ctmp_sva_1[38:0]),
          attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_38_0, GEMM_3D_FLOAT_LOOP_3_1_and_52_nl,
          attention_2_1_16_16_4_4_attn_output_0_0_3_sva_2_mx1_38_0, {apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c0
          , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_lpi_3_mx0c1 , for_for_and_22_nl
          , and_dcpl_548 , and_dcpl_207 , and_dcpl_220 , and_dcpl_222 , and_dcpl_187});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_attn_output_and_25_cse ) begin
      attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3 <= MUX1HOT_v_40_7_2(({{10{strm_in_rsci_idat_mxwt[29]}},
          strm_in_rsci_idat_mxwt}), input_0_1_sva_1, attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1,
          attention_2_1_16_16_4_4_k_embed_1_0_2_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2,
          GEMM_3D_FLOAT_LOOP_3_1_and_28_nl, attention_2_1_16_16_4_4_attn_output_1_0_3_sva_2_mx1,
          {and_521_nl , and_523_nl , and_dcpl_346 , and_dcpl_204 , and_dcpl_220 ,
          and_dcpl_222 , and_dcpl_187});
      attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3 <= MUX1HOT_v_40_7_2(({{10{strm_in_rsci_idat_mxwt[29]}},
          strm_in_rsci_idat_mxwt}), input_0_14_sva_1, attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1,
          attention_2_1_16_16_4_4_k_embed_1_0_3_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2,
          GEMM_3D_FLOAT_LOOP_3_1_and_29_nl, attention_2_1_16_16_4_4_attn_output_2_0_0_sva_2_mx1,
          {and_527_nl , and_529_nl , and_dcpl_346 , and_dcpl_204 , and_dcpl_220 ,
          and_dcpl_222 , and_dcpl_187});
      attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3 <= MUX1HOT_v_40_7_2(({{10{strm_in_rsci_idat_mxwt[29]}},
          strm_in_rsci_idat_mxwt}), input_0_6_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1,
          attention_2_1_16_16_4_4_k_embed_2_0_0_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2,
          GEMM_3D_FLOAT_LOOP_3_1_and_31_nl, attention_2_1_16_16_4_4_attn_output_2_0_1_sva_2_mx1,
          {and_531_nl , and_533_nl , and_dcpl_346 , and_dcpl_204 , and_dcpl_220 ,
          and_dcpl_222 , and_dcpl_187});
      attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3 <= MUX1HOT_v_40_7_2(({{10{strm_in_rsci_idat_mxwt[29]}},
          strm_in_rsci_idat_mxwt}), input_0_9_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1,
          attention_2_1_16_16_4_4_k_embed_2_0_1_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2,
          GEMM_3D_FLOAT_LOOP_3_1_and_33_nl, attention_2_1_16_16_4_4_attn_output_2_0_2_sva_2_mx1,
          {and_535_nl , and_537_nl , and_dcpl_346 , and_dcpl_204 , and_dcpl_220 ,
          and_dcpl_222 , and_dcpl_187});
      attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3 <= MUX1HOT_v_40_7_2(({{10{strm_in_rsci_idat_mxwt[29]}},
          strm_in_rsci_idat_mxwt}), input_0_5_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1,
          attention_2_1_16_16_4_4_k_embed_2_0_2_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2,
          GEMM_3D_FLOAT_LOOP_3_1_and_35_nl, attention_2_1_16_16_4_4_attn_output_2_0_3_sva_2_mx1,
          {and_539_nl , and_541_nl , and_dcpl_346 , and_dcpl_204 , and_dcpl_220 ,
          and_dcpl_222 , and_dcpl_187});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_995)
        | attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c0 | attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c1
        | and_dcpl_346 | and_dcpl_204 | attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c5
        | and_dcpl_222 | and_dcpl_187 | attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c8
        | attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c10) & mux_1133_nl )
        begin
      attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          mux_nl, nor_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_997)
        | attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c0 | attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c1
        | and_dcpl_346 | (~ mux_1147_itm) | and_dcpl_204 | and_dcpl_524 | and_dcpl_222
        | and_dcpl_187 | mux_tmp_1163 | attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c10)
        ) begin
      attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          mux1h_nl, not_4622_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_999)
        | attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c0 | attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c1
        | and_dcpl_346 | (~ mux_1177_itm) | and_dcpl_204 | and_dcpl_524 | and_dcpl_222
        | and_dcpl_187 | mux_tmp_1163 | attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c10)
        ) begin
      attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          mux1h_1_nl, not_4624_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_1000)
        | attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c0 | attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c1
        | and_dcpl_242 | (~ mux_1197_itm) | and_dcpl_344 | and_dcpl_346 | and_dcpl_204
        | and_dcpl_524 | and_dcpl_222 | and_dcpl_187 | attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c10
        | attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c12) ) begin
      attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          mux1h_2_nl, not_4626_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4 <= 1'b0;
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0 <= 4'b0000;
    end
    else if ( LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_1_ssc ) begin
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4 <= (LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_7_nl
          & (~ and_dcpl_477) & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_nand_seb) | and_585_seb;
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0 <= MUX_v_4_2_2(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_4_nl,
          4'b1111, and_585_seb);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1 <= 5'b00000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (and_dcpl_415 |
        and_dcpl_257) ) begin
      LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1 <= MUX_v_5_2_2(LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp,
          RMS_NORM_LOOP_2_2_acc_1_tmp, and_dcpl_257);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_abs_qr_35_0_lpi_1_dfm_35 <= 1'b0;
      attention_abs_qr_35_0_lpi_1_dfm_34_0 <= 35'b00000000000000000000000000000000000;
    end
    else if ( attention_abs_qelse_and_ssc ) begin
      attention_abs_qr_35_0_lpi_1_dfm_35 <= (attention_abs_qr_35_0_lpi_1_dfm_mx0w0[35])
          & (~ attention_abs_qr_35_0_lpi_1_dfm_mx0c1);
      attention_abs_qr_35_0_lpi_1_dfm_34_0 <= MUX_v_35_2_2((attention_abs_qr_35_0_lpi_1_dfm_mx0w0[34:0]),
          (operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1[34:0]),
          attention_abs_qr_35_0_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      compute_sqrt_guess_sva_34 <= 1'b0;
      compute_sqrt_guess_sva_33_0 <= 34'b0000000000000000000000000000000000;
    end
    else if ( compute_sqrt_guess_and_ssc ) begin
      compute_sqrt_guess_sva_34 <= MUX_s_1_2_2(attention_abs_qr_35_0_lpi_1_dfm_mx1_35,
          (compute_sqrt_for_acc_1_itm_40_1_1[34]), and_dcpl_290);
      compute_sqrt_guess_sva_33_0 <= MUX_v_34_2_2(attention_abs_qr_35_0_lpi_1_dfm_mx1_34_1,
          (compute_sqrt_for_acc_1_itm_40_1_1[33:0]), and_dcpl_290);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_15
          <= 1'b0;
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd
          <= 3'b000;
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1
          <= 3'b000;
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2
          <= 1'b0;
    end
    else if ( operator_40_24_true_AC_TRN_AC_WRAP_1_and_ssc ) begin
      operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_15
          <= MUX_s_1_2_2((operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z[15]), attention_2_1_16_16_4_4_q_proj_attention_2_1_16_16_4_4_q_proj_mux_12_nl,
          and_622_rgt);
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd
          <= MUX1HOT_v_3_4_2((operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z[14:12]),
          attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_14_12, (z_out[14:12]), (APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_itm[14:12]),
          {and_615_itm , operator_40_24_true_AC_TRN_AC_WRAP_1_and_4_cse , and_1191_rgt
          , and_dcpl_583});
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1
          <= MUX1HOT_v_3_5_2((operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z[11:9]),
          (operator_40_24_true_AC_TRN_AC_WRAP_1_conc_1_itm_11_0[11:9]), attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_11_9,
          (z_out[11:9]), (APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_itm[11:9]),
          {and_615_itm , and_dcpl_438 , operator_40_24_true_AC_TRN_AC_WRAP_1_and_4_cse
          , and_1191_rgt , and_dcpl_583});
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2
          <= MUX1HOT_s_1_6_2((operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z[8]),
          (operator_40_24_true_AC_TRN_AC_WRAP_1_conc_1_itm_11_0[8]), attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_8,
          (z_out[8]), (APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_itm[8]),
          (operator_40_24_true_AC_TRN_AC_WRAP_1_conc_3_itm_8_0[8]), {and_615_itm
          , and_dcpl_438 , operator_40_24_true_AC_TRN_AC_WRAP_1_and_4_cse , and_1191_rgt
          , and_dcpl_583 , and_dcpl_448});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3
          <= 8'b00000000;
    end
    else if ( operator_40_24_true_AC_TRN_AC_WRAP_1_and_ssc & (~((~ mux_1309_cse)
        & and_dcpl_383 & and_dcpl_338 & and_dcpl_576)) ) begin
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3
          <= MUX1HOT_v_8_8_2((operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z[7:0]),
          (operator_40_24_true_AC_TRN_AC_WRAP_1_conc_1_itm_11_0[7:0]), LINEAR_FORWARD_NO_MUL_LOOP_3_1_packed_val_read_rom_k_weights_rom_map_1_itm,
          LINEAR_FORWARD_NO_MUL_LOOP_3_3_packed_val_read_rom_o_weights_rom_map_1_itm,
          attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0, (z_out[7:0]), (APPLY_ROTARY_POS_EMB_LOOP_6_cosval_read_rom_cos_tab_rom_map_1_itm[7:0]),
          (operator_40_24_true_AC_TRN_AC_WRAP_1_conc_3_itm_8_0[7:0]), {and_615_itm
          , and_dcpl_438 , operator_40_24_true_AC_TRN_AC_WRAP_1_and_2_nl , and_dcpl_739
          , operator_40_24_true_AC_TRN_AC_WRAP_1_and_4_cse , and_1191_rgt , and_dcpl_583
          , and_dcpl_448});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_38_0 <= 39'b000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & and_dcpl_344 )
        begin
      QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_38_0 <= QUANTIZE_ACTIVATION_LOOP_1_max_val_lpi_2_dfm_1_38_0_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_quantized_hidden_states_0_9_sva_7 <= 1'b0;
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_hidden_states_and_ssc ) begin
      attention_2_1_16_16_4_4_quantized_hidden_states_0_9_sva_7 <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_cse;
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_9_1_cse <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_quantized_hidden_states_0_6_sva_7 <= 1'b0;
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_hidden_states_and_1_ssc ) begin
      attention_2_1_16_16_4_4_quantized_hidden_states_0_6_sva_7 <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_cse;
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_6_1_cse <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_quantized_hidden_states_0_8_sva_7 <= 1'b0;
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_hidden_states_and_2_ssc ) begin
      attention_2_1_16_16_4_4_quantized_hidden_states_0_8_sva_7 <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_cse;
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_8_1_cse <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_quantized_hidden_states_0_7_sva_7 <= 1'b0;
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_hidden_states_and_3_ssc ) begin
      attention_2_1_16_16_4_4_quantized_hidden_states_0_7_sva_7 <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_cse;
      reg_attention_2_1_16_16_4_4_quantized_hidden_states_0_7_1_cse <= INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd <= 3'b000;
    end
    else if ( RMS_NORM_LOOP_2_2_i_and_ssc ) begin
      reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd <= MUX_v_3_2_2(3'b000, RMS_NORM_LOOP_2_2_i_mux1h_3_nl,
          RMS_NORM_LOOP_2_2_i_not_2_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 <= 1'b0;
    end
    else if ( RMS_NORM_LOOP_2_2_i_and_ssc & (~(and_dcpl_1151 | ((~ and_dcpl_557)
        & RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c4))) ) begin
      reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 <= RMS_NORM_LOOP_2_2_i_mux1h_6_nl
          & (~ RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      RMS_NORM_LOOP_2_2_i_4_0_sva_1 <= 5'b00000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1434_nl |
        (fsm_output[8])) ) begin
      RMS_NORM_LOOP_2_2_i_4_0_sva_1 <= MUX_v_5_2_2(RMS_NORM_LOOP_2_2_acc_1_tmp, LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp,
          and_dcpl_257);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1 <= 1'b0;
      reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 <= 1'b0;
    end
    else if ( CACHE_UPDATE_LOOP_3_k_and_ssc ) begin
      reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1_1 <= MUX1HOT_s_1_3_2((z_out_3[2]), (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3[2]),
          (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[2]), {and_dcpl_318 , and_dcpl_328 , and_dcpl_635});
      reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 <= MUX1HOT_s_1_4_2(QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_3_nl,
          (z_out_3[1]), (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3[1]), (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[1]),
          {CACHE_UPDATE_LOOP_3_k_2_0_sva_1_mx0c1 , and_dcpl_318 , and_dcpl_328 ,
          and_dcpl_635});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 <= 1'b0;
    end
    else if ( CACHE_UPDATE_LOOP_3_k_and_ssc & (~(and_dcpl_629 | compute_sqrt_for_i_and_2_cse))
        ) begin
      reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1 <= MUX1HOT_s_1_6_2(RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_and_nl,
          QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_4_nl, (z_out_3[0]),
          (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_14_sdt_mx0w3[0]), (GEMM_3D_FLOAT_LOOP_3_acc_6_tmp[0]),
          (~ QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1),
          {CACHE_UPDATE_LOOP_3_k_and_1_nl , CACHE_UPDATE_LOOP_3_k_2_0_sva_1_mx0c1
          , and_dcpl_318 , and_dcpl_328 , and_dcpl_635 , and_dcpl_557});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd <= 1'b0;
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 <= 1'b0;
    end
    else if ( GEMM_3D_FLOAT_LOOP_1_i_and_ssc ) begin
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd <= (z_out_5[1]) & (~ GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c2);
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 <= GEMM_3D_FLOAT_LOOP_1_i_mux_1_nl
          & (~ GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c2);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_0_0_sva_2 <= 40'b0000000000000000000000000000000000000000;
      input_0_1_sva_2 <= 40'b0000000000000000000000000000000000000000;
      input_0_2_sva_2_39 <= 1'b0;
      input_0_2_sva_2_38_0 <= 39'b000000000000000000000000000000000000000;
      input_0_3_sva_2 <= 40'b0000000000000000000000000000000000000000;
      input_0_4_sva_2 <= 40'b0000000000000000000000000000000000000000;
      input_0_5_sva_2 <= 40'b0000000000000000000000000000000000000000;
      input_0_6_sva_2 <= 40'b0000000000000000000000000000000000000000;
      input_0_7_sva_2 <= 40'b0000000000000000000000000000000000000000;
      input_0_8_sva_2 <= 40'b0000000000000000000000000000000000000000;
      input_0_9_sva_2 <= 40'b0000000000000000000000000000000000000000;
      input_0_10_sva_2 <= 40'b0000000000000000000000000000000000000000;
      input_0_11_sva_2 <= 40'b0000000000000000000000000000000000000000;
      input_0_12_sva_2 <= 40'b0000000000000000000000000000000000000000;
      input_0_13_sva_2_39 <= 1'b0;
      input_0_13_sva_2_38_0 <= 39'b000000000000000000000000000000000000000;
      input_0_14_sva_2 <= 40'b0000000000000000000000000000000000000000;
      input_0_15_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( input_and_28_cse ) begin
      input_0_0_sva_2 <= MUX_v_40_2_2((z_out_13_71_28[39:0]), attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1,
          and_688_nl);
      input_0_1_sva_2 <= MUX_v_40_2_2((z_out_13_71_28[39:0]), input_0_1_sva_1, and_693_nl);
      input_0_2_sva_2_39 <= MUX_s_1_2_2((z_out_13_71_28[39]), input_0_2_sva_1_39,
          and_699_ssc);
      input_0_2_sva_2_38_0 <= MUX_v_39_2_2((z_out_13_71_28[38:0]), input_0_2_sva_1_38_0,
          and_699_ssc);
      input_0_3_sva_2 <= MUX_v_40_2_2((z_out_13_71_28[39:0]), input_0_3_sva_1, and_704_nl);
      input_0_4_sva_2 <= MUX_v_40_2_2((z_out_13_71_28[39:0]), input_0_4_sva_1, and_709_nl);
      input_0_5_sva_2 <= MUX_v_40_2_2((z_out_13_71_28[39:0]), input_0_5_sva_1, and_713_nl);
      input_0_6_sva_2 <= MUX_v_40_2_2((z_out_13_71_28[39:0]), input_0_6_sva_1, and_717_nl);
      input_0_7_sva_2 <= MUX_v_40_2_2((z_out_13_71_28[39:0]), input_0_7_sva_1, and_721_nl);
      input_0_8_sva_2 <= MUX_v_40_2_2((z_out_13_71_28[39:0]), input_0_8_sva_1, and_725_nl);
      input_0_9_sva_2 <= MUX_v_40_2_2((z_out_13_71_28[39:0]), input_0_9_sva_1, and_729_nl);
      input_0_10_sva_2 <= MUX_v_40_2_2((z_out_13_71_28[39:0]), input_0_10_sva_1,
          and_733_nl);
      input_0_11_sva_2 <= MUX_v_40_2_2((z_out_13_71_28[39:0]), input_0_11_sva_1,
          and_737_nl);
      input_0_12_sva_2 <= MUX_v_40_2_2((z_out_13_71_28[39:0]), input_0_12_sva_1,
          and_741_nl);
      input_0_13_sva_2_39 <= MUX_s_1_2_2((z_out_13_71_28[39]), input_0_13_sva_1_39,
          and_745_ssc);
      input_0_13_sva_2_38_0 <= MUX_v_39_2_2((z_out_13_71_28[38:0]), input_0_13_sva_1_38_0,
          and_745_ssc);
      input_0_14_sva_2 <= MUX_v_40_2_2((z_out_13_71_28[39:0]), input_0_14_sva_1,
          and_749_nl);
      input_0_15_sva_1 <= MUX_v_40_2_2((z_out_13_71_28[39:0]), attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3,
          and_753_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~(or_tmp_833 |
        nand_197_cse | or_dcpl_1109 | or_1984_cse)) ) begin
      RMS_NORM_LOOP_2_slc_RMS_NORM_LOOP_2_mul_67_28_ncse_sva <= z_out_13_71_28[39:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 <= 1'b0;
    end
    else if ( APPLY_ROTARY_POS_EMB_LOOP_1_i_and_ssc ) begin
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd <= (z_out_4[1]) & mux_1512_itm;
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 <= APPLY_ROTARY_POS_EMB_LOOP_1_i_mux1h_5_nl
          & mux_1512_itm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd <= 1'b0;
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_1 <= 1'b0;
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_2 <= 1'b0;
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_3 <= 1'b0;
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_4 <= 1'b0;
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_5 <= 1'b0;
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_6 <= 1'b0;
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_q_proj_and_4_ssc ) begin
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1,
          attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_7,
          {nor_1144_itm , and_dcpl_240 , and_dcpl_626});
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_1 <= MUX1HOT_s_1_3_2((~
          QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_6,
          attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_6, {nor_1144_itm , and_dcpl_240
          , and_dcpl_626});
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_2 <= MUX1HOT_s_1_3_2((~
          QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_5,
          attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_5, {nor_1144_itm , and_dcpl_240
          , and_dcpl_626});
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_3 <= MUX1HOT_s_1_3_2((~
          QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_4,
          attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_4, {nor_1144_itm , and_dcpl_240
          , and_dcpl_626});
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_4 <= MUX1HOT_s_1_3_2((~
          QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_3,
          attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_3, {nor_1144_itm , and_dcpl_240
          , and_dcpl_626});
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_5 <= MUX1HOT_s_1_3_2((~
          QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_2,
          attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_2, {nor_1144_itm , and_dcpl_240
          , and_dcpl_626});
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_6 <= MUX1HOT_s_1_3_2((~
          QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_1,
          attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_1, {nor_1144_itm , and_dcpl_240
          , and_dcpl_626});
      reg_attention_2_1_16_16_4_4_q_proj_1_0_0_lpi_3_15_0_1_ftd_7 <= MUX1HOT_s_1_3_2((~
          QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_0_mx0w1_0,
          attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_0, {nor_1144_itm , and_dcpl_240
          , and_dcpl_626});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_v_proj_re_and_cse ) begin
      attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_4_nl, not_4557_nl);
      attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_8_nl, not_4558_nl);
      attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_12_nl, not_4559_nl);
      attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_16_nl, not_4560_nl);
      attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_20_nl, not_4561_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_21_nl, not_4562_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_3_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_q_proj_re_and_cse ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_35_nl, not_4441_nl);
      attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_34_nl, not_4440_nl);
      attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_33_nl, not_4439_nl);
      attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_32_nl, not_4438_nl);
      attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_31_nl, not_4437_nl);
      attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_30_nl, not_4436_nl);
      attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_29_nl, not_4435_nl);
      attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_28_nl, not_4434_nl);
      attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_27_nl, not_4433_nl);
      attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_26_nl, not_4432_nl);
      attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_25_nl, not_4431_nl);
      attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_24_nl, not_4430_nl);
      attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_23_nl, not_4429_nl);
      attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_22_nl, not_4428_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_3_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_7_sva_2_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_proj_re_and_1_cse ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_21_nl, not_4427_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_20_nl, not_4426_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_19_nl, not_4425_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_18_nl, not_4424_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_17_nl, not_4422_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux_16_nl, not_4415_nl);
      attention_2_1_16_16_4_4_k_proj_re_0_7_sva_2_39_16 <= MUX_v_24_2_2((rms_norm_16_div_cmp_z_oreg[39:16]),
          attention_2_1_16_16_4_4_k_proj_re_0_7_sva_1_39_16, and_1184_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (and_dcpl_619 |
        attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16_mx0c1 | and_dcpl_843 |
        and_dcpl_207 | and_dcpl_847) ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_40_nl, not_4423_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (and_dcpl_619 |
        attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16_mx0c1 | and_dcpl_856 |
        and_dcpl_207 | and_dcpl_847) ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_42_nl, not_4421_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (and_dcpl_619 |
        attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16_mx0c1 | and_dcpl_860 |
        and_dcpl_207 | and_dcpl_847) ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_43_nl, not_4420_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (and_dcpl_619 |
        attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16_mx0c1 | and_dcpl_864 |
        and_dcpl_207 | and_dcpl_847) ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_44_nl, not_4419_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (and_dcpl_619 |
        attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16_mx0c1 | and_dcpl_868 |
        and_dcpl_207 | and_dcpl_847) ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_45_nl, not_4418_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (and_dcpl_619 |
        attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16_mx0c1 | and_dcpl_872 |
        and_dcpl_207 | and_dcpl_847) ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_46_nl, not_4417_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (and_dcpl_619 |
        attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16_mx0c1 | and_dcpl_876 |
        and_dcpl_207 | and_dcpl_847) ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_47_nl, not_4416_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 <= 1'b0;
    end
    else if ( APPLY_ROTARY_POS_EMB_LOOP_6_k_and_ssc ) begin
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd <= GEMM_3D_FLOAT_LOOP_4_l_GEMM_3D_FLOAT_LOOP_4_l_mux_nl
          & (~ APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c0);
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 <= GEMM_3D_FLOAT_LOOP_4_l_mux1h_13_nl
          & (~ APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c0);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1641_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_26_nl, not_4471_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1644_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_28_nl, not_4470_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1727_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_40_nl, not_4464_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1816_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_43_nl, not_4458_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1825_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_42_nl, not_4457_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1834_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_41_nl, not_4456_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1843_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_40_nl, not_4455_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1852_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_39_nl, not_4454_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1861_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_38_nl, not_4453_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1870_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_37_nl, not_4452_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1878_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_36_nl, not_4451_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1887_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_35_nl, not_4450_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1896_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_34_nl, not_4449_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1905_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_33_nl, not_4448_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1914_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_32_nl, not_4447_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1923_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_31_nl, not_4446_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1932_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_30_nl, not_4445_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_1941_nl |
        (fsm_output[8])) ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux_29_nl, not_4444_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~((~ mux_1946_nl)
        & and_dcpl_259)) ) begin
      attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_66_nl, not_4563_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~((~ mux_1947_nl)
        & and_dcpl_259)) ) begin
      attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_67_nl, not_4564_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_1068)
        | and_dcpl_619 | apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c1
        | and_dcpl_983 | and_dcpl_240 | and_dcpl_626 | and_dcpl_739 | apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c8)
        & (~ mux_1973_nl) ) begin
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          ({attention_2_1_16_16_4_4_k_proj_re_mux1h_69_nl , attention_2_1_16_16_4_4_k_proj_re_mux1h_119_nl}),
          not_4565_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_15_8 <= 8'b00000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_7 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_6 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_5 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_4 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_3 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_2 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_1 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_0 <= 1'b0;
    end
    else if ( apply_rotary_pos_emb_1_4_4_rotated_q_and_16_ssc ) begin
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_15_8 <= MUX_v_8_2_2(8'b00000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_70_nl, not_5074_nl);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_7 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_128_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_6 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_129_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_5 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_130_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_4 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_131_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_3 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_132_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_2 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_133_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_1 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_134_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_0 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_135_nl
          & (~ and_dcpl_619);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_8 <= 8'b00000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_7 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_6 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_5 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_4 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_3 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_2 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_1 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_0 <= 1'b0;
    end
    else if ( apply_rotary_pos_emb_1_4_4_rotated_q_and_17_ssc ) begin
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_8 <= MUX_v_8_2_2(8'b00000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_71_nl, not_5066_nl);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_7 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_120_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_6 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_121_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_5 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_122_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_4 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_123_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_3 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_124_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_2 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_125_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_1 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_126_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_0 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_127_nl
          & (~ and_dcpl_619);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_1145)
        | and_dcpl_619 | attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c1 |
        and_dcpl_410 | and_dcpl_739 | attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c6)
        & mux_2012_nl ) begin
      attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_72_nl, not_4566_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~(or_dcpl_1146
        | (~(mux_2022_nl | (fsm_output[8]))))) | and_dcpl_619 | attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0_mx0c1
        | and_dcpl_410) ) begin
      attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_73_nl, not_4567_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8 <= 8'b00000000;
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7 <= 1'b0;
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6 <= 1'b0;
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5 <= 1'b0;
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4 <= 1'b0;
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3 <= 1'b0;
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2 <= 1'b0;
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1 <= 1'b0;
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0 <= 1'b0;
    end
    else if ( APPLY_ROTARY_POS_EMB_LOOP_6_and_30_ssc ) begin
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8 <= MUX_v_8_2_2(8'b00000000, attention_2_1_16_16_4_4_k_proj_re_mux1h_74_nl,
          not_5054_nl);
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_117_nl
          & (~ and_dcpl_619);
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_152_nl
          & (~ and_dcpl_619);
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_153_nl
          & (~ and_dcpl_619);
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_154_nl
          & (~ and_dcpl_619);
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_155_nl
          & (~ and_dcpl_619);
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_156_nl
          & (~ and_dcpl_619);
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_157_nl
          & (~ and_dcpl_619);
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_158_nl
          & (~ and_dcpl_619);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd <= 3'b000;
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1 <= 13'b0000000000000;
    end
    else if ( apply_rotary_pos_emb_1_4_4_rotated_q_and_18_ssc ) begin
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd <= MUX_v_3_2_2(3'b000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_75_nl, not_4569_nl);
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1 <= MUX_v_13_2_2(13'b0000000000000,
          ({attention_2_1_16_16_4_4_k_proj_re_mux1h_116_nl , attention_2_1_16_16_4_4_k_proj_re_mux1h_144_nl
          , attention_2_1_16_16_4_4_k_proj_re_mux1h_145_nl , attention_2_1_16_16_4_4_k_proj_re_mux1h_146_nl
          , attention_2_1_16_16_4_4_k_proj_re_mux1h_147_nl , attention_2_1_16_16_4_4_k_proj_re_mux1h_148_nl
          , attention_2_1_16_16_4_4_k_proj_re_mux1h_149_nl , attention_2_1_16_16_4_4_k_proj_re_mux1h_150_nl
          , attention_2_1_16_16_4_4_k_proj_re_mux1h_151_nl}), not_5062_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_15_8 <= 8'b00000000;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_7 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_6 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_5 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_4 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_3 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_2 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_1 <= 1'b0;
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_0 <= 1'b0;
    end
    else if ( apply_rotary_pos_emb_1_4_4_rotated_q_and_19_ssc ) begin
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_15_8 <= MUX_v_8_2_2(8'b00000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_76_nl, not_5088_nl);
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_7 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_136_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_6 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_137_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_5 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_138_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_4 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_139_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_3 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_140_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_2 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_141_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_1 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_142_nl
          & (~ and_dcpl_619);
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_0 <= attention_2_1_16_16_4_4_k_proj_re_mux1h_143_nl
          & (~ and_dcpl_619);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~((~ mux_2038_nl)
        & and_dcpl_259)) ) begin
      attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_77_nl, not_4571_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~((~ mux_2039_nl)
        & and_dcpl_259)) ) begin
      attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_78_nl, not_4572_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~((~ mux_2040_nl)
        & and_dcpl_259)) ) begin
      attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_79_nl, not_4573_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_2051_nl |
        (fsm_output[7])) ) begin
      attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_80_nl, not_4574_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~((~ mux_2052_nl)
        & and_dcpl_259)) ) begin
      attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_81_nl, not_4575_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~((~ mux_2053_nl)
        & and_dcpl_259)) ) begin
      attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_82_nl, not_4576_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~((~ mux_2054_nl)
        & and_dcpl_259)) ) begin
      attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_83_nl, not_4577_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~((~ mux_2055_nl)
        & and_dcpl_259)) ) begin
      attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_15_0 <= MUX_v_16_2_2(16'b0000000000000000,
          attention_2_1_16_16_4_4_k_proj_re_mux1h_84_nl, not_4578_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (mux_2059_nl |
        (fsm_output[8])) ) begin
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_51_nl, not_4414_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~(or_dcpl_1068
        | (~(mux_2063_nl | (fsm_output[8]))))) | and_dcpl_619 | apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16_mx0c1
        | and_dcpl_1003) ) begin
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_52_nl, not_4413_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~((~ mux_2068_nl)
        & and_dcpl_581)) ) begin
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_53_nl, not_4412_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~(or_dcpl_1068
        | ((~ mux_tmp_2067) & and_dcpl_581))) | and_dcpl_619 | apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16_mx0c1
        | and_dcpl_959) ) begin
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_54_nl, not_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~(or_dcpl_1145
        | and_dcpl_1055)) | and_dcpl_619 | and_dcpl_726 | and_dcpl_410) ) begin
      attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_55_nl, not_4579_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (and_dcpl_619 |
        and_dcpl_726 | and_dcpl_257 | and_dcpl_1033 | and_dcpl_983 | and_dcpl_240
        | and_dcpl_1034 | and_dcpl_207 | and_dcpl_213 | and_dcpl_583 | and_dcpl_265)
        ) begin
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_56_nl, not_4580_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (and_dcpl_619 |
        and_dcpl_726 | and_dcpl_257 | and_dcpl_1011 | and_dcpl_983 | and_dcpl_240
        | and_dcpl_207 | and_dcpl_847 | and_dcpl_583) ) begin
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16 <= MUX_v_24_2_2(24'b000000000000000000000000,
          attention_2_1_16_16_4_4_v_proj_re_mux1h_57_nl, not_4581_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_7 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_6 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_5 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_4 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_3 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_2 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_1 <= 1'b0;
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_0 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_q_proj_and_5_ssc ) begin
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_7 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_nl,
          attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_7, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_7,
          {nor_1228_ssc , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_6 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse,
          attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_6, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_6,
          {nor_1228_ssc , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_5 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse,
          attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_5, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_5,
          {nor_1228_ssc , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_4 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse,
          attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_4, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_4,
          {nor_1228_ssc , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_3 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse,
          attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_3, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_3,
          {nor_1228_ssc , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_2 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse,
          attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_2, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_2,
          {nor_1228_ssc , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_1 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse,
          attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_1, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_1,
          {nor_1228_ssc , and_dcpl_240 , and_dcpl_626});
      attention_2_1_16_16_4_4_q_proj_2_0_3_lpi_3_0 <= MUX1HOT_s_1_3_2(QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_1_cse,
          attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_0_mx0w1_0, attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_0,
          {nor_1228_ssc , and_dcpl_240 , and_dcpl_626});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd <= 8'b00000000;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd <= 8'b00000000;
    end
    else if ( APPLY_ROTARY_POS_EMB_LOOP_6_and_28_cse ) begin
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd <= MUX1HOT_v_8_6_2((drf_output_sdt_2_sva_15_0_mx0w0[15:8]),
          attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_8, attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_15_8,
          apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8,
          apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_8, APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_nl,
          {and_dcpl_257 , and_dcpl_1073 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847
          , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd <= MUX1HOT_v_8_6_2((z_out[15:8]),
          attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_8, attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_15_8,
          apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8,
          apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_8, APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_nl,
          {and_dcpl_257 , and_dcpl_1073 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847
          , and_dcpl_583});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1 <= 1'b0;
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0 <= 1'b0;
    end
    else if ( APPLY_ROTARY_POS_EMB_LOOP_6_and_31_cse ) begin
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm[7]),
          (drf_output_sdt_2_sva_15_0_mx0w0[7]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_7,
          attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_7, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7,
          apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_7, APPLY_ROTARY_POS_EMB_LOOP_6_mux_66_nl,
          {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073 , and_dcpl_240 , and_dcpl_207
          , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm[6]),
          (drf_output_sdt_2_sva_15_0_mx0w0[6]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_6,
          attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_6, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6,
          apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_6, APPLY_ROTARY_POS_EMB_LOOP_6_mux_74_nl,
          {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073 , and_dcpl_240 , and_dcpl_207
          , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm[5]),
          (drf_output_sdt_2_sva_15_0_mx0w0[5]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_5,
          attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_5, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5,
          apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_5, APPLY_ROTARY_POS_EMB_LOOP_6_mux_75_nl,
          {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073 , and_dcpl_240 , and_dcpl_207
          , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm[4]),
          (drf_output_sdt_2_sva_15_0_mx0w0[4]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_4,
          attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_4, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4,
          apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_4, APPLY_ROTARY_POS_EMB_LOOP_6_mux_76_nl,
          {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073 , and_dcpl_240 , and_dcpl_207
          , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm[3]),
          (drf_output_sdt_2_sva_15_0_mx0w0[3]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_3,
          attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_3, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3,
          apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_3, APPLY_ROTARY_POS_EMB_LOOP_6_mux_77_nl,
          {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073 , and_dcpl_240 , and_dcpl_207
          , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm[2]),
          (drf_output_sdt_2_sva_15_0_mx0w0[2]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_2,
          attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_2, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2,
          apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_2, APPLY_ROTARY_POS_EMB_LOOP_6_mux_78_nl,
          {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073 , and_dcpl_240 , and_dcpl_207
          , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm[1]),
          (drf_output_sdt_2_sva_15_0_mx0w0[1]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_1,
          attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_1, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1,
          apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_1, APPLY_ROTARY_POS_EMB_LOOP_6_mux_79_nl,
          {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073 , and_dcpl_240 , and_dcpl_207
          , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_2_packed_val_read_rom_v_weights_rom_map_1_itm[0]),
          (drf_output_sdt_2_sva_15_0_mx0w0[0]), attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_0,
          attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_0_mx0w1_0, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0,
          apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_0, APPLY_ROTARY_POS_EMB_LOOP_6_mux_80_nl,
          {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073 , and_dcpl_240 , and_dcpl_207
          , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm[7]),
          (z_out[7]), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd,
          attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_7, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7,
          reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_61_nl, {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073
          , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm[6]),
          (z_out[6]), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_1,
          attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_6, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6,
          reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_1,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_81_nl, {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073
          , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm[5]),
          (z_out[5]), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_2,
          attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_5, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5,
          reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_2,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_82_nl, {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073
          , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm[4]),
          (z_out[4]), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_3,
          attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_4, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4,
          reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_3,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_83_nl, {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073
          , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm[3]),
          (z_out[3]), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_4,
          attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_3, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3,
          reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_4,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_84_nl, {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073
          , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm[2]),
          (z_out[2]), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_5,
          attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_2, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2,
          reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_5,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_85_nl, {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073
          , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm[1]),
          (z_out[1]), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_6,
          attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_1, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1,
          reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_6,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_86_nl, {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073
          , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583});
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0 <= MUX1HOT_s_1_7_2((LINEAR_FORWARD_NO_MUL_LOOP_3_packed_val_read_rom_q_weights_rom_map_1_itm[0]),
          (z_out[0]), reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_7,
          attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_mx0w1_0, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0,
          reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_7,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_87_nl, {and_dcpl_888 , and_dcpl_257 , and_dcpl_1073
          , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_0_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_14_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_13_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_12_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_11_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_4_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_10_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_5_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_9_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_6_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_8_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_7_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_q_proj_re_0_15_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_q_proj_re_and_29_cse ) begin
      attention_2_1_16_16_4_4_q_proj_re_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_14_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_13_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_2_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_12_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_11_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_4_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_10_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_5_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_9_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_6_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_8_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_7_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_q_proj_re_0_15_sva_1_39_16 <= attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_39_16_mx1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_15_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_0_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_14_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_13_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_12_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_11_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_4_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_10_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_5_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_9_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_6_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_8_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_k_proj_re_0_7_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_proj_re_and_65_cse ) begin
      attention_2_1_16_16_4_4_k_proj_re_0_15_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_14_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_13_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_2_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_12_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_3_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_11_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_4_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_10_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_5_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_9_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_6_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_8_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_k_proj_re_0_7_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16_mx1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_v_proj_re_0_15_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_0_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_14_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_13_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_12_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_4_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_10_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_5_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_9_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_6_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_8_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_7_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_v_proj_re_and_32_cse ) begin
      attention_2_1_16_16_4_4_v_proj_re_0_15_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_14_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_14_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_13_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_13_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_2_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_2_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_12_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_12_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_3_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_11_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_4_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_4_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_10_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_10_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_5_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_5_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_9_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_6_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_6_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_8_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_39_16_mx1;
      attention_2_1_16_16_4_4_v_proj_re_0_7_sva_1_39_16 <= attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16_mx1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      LINEAR_FORWARD_NO_MUL_LOOP_2_mul_itm <= 60'b000000000000000000000000000000000000000000000000000000000000;
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_mul_mut <= 60'b000000000000000000000000000000000000000000000000000000000000;
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut <= 61'b0000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( LINEAR_FORWARD_NO_MUL_LOOP_2_and_cse ) begin
      LINEAR_FORWARD_NO_MUL_LOOP_2_mul_itm <= z_out_10[59:0];
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_mul_mut <= z_out_9;
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut <= LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8 <= 8'b00000000;
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd <= 1'b0;
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1 <= 1'b0;
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2 <= 1'b0;
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3 <= 1'b0;
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4 <= 1'b0;
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5 <= 1'b0;
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6 <= 1'b0;
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7 <= 1'b0;
    end
    else if ( LINEAR_FORWARD_NO_MUL_LOOP_2_1_and_29_ssc ) begin
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8 <= MUX1HOT_v_8_7_2((z_out_1[15:8]),
          attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_15_8, RESHAPE_2D_TO_3D_LOOP_3_1_mux_13_cse,
          apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_8, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8,
          ({APPLY_ROTARY_POS_EMB_LOOP_6_mux_32_nl , APPLY_ROTARY_POS_EMB_LOOP_6_mux_70_nl
          , APPLY_ROTARY_POS_EMB_LOOP_6_mux_71_nl , APPLY_ROTARY_POS_EMB_LOOP_6_mux_72_nl}),
          (drf_output_sdt_3_sva_15_0_mx0w3[15:8]), {and_dcpl_257 , operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse
          , and_dcpl_240 , attention_2_1_16_16_4_4_k_proj_re_or_17_cse , and_dcpl_207
          , and_dcpl_583 , and_dcpl_265});
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd <= MUX1HOT_s_1_7_2((z_out_1[7]),
          attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_7, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_7,
          apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_7, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_7,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_50_nl, (drf_output_sdt_3_sva_15_0_mx0w3[7]),
          {and_dcpl_257 , operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse ,
          and_dcpl_240 , attention_2_1_16_16_4_4_k_proj_re_or_17_cse , and_dcpl_207
          , and_dcpl_583 , and_dcpl_265});
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1 <= MUX1HOT_s_1_7_2((z_out_1[6]),
          attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_6, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_6,
          apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_6, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_6,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_51_nl, (drf_output_sdt_3_sva_15_0_mx0w3[6]),
          {and_dcpl_257 , operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse ,
          and_dcpl_240 , attention_2_1_16_16_4_4_k_proj_re_or_17_cse , and_dcpl_207
          , and_dcpl_583 , and_dcpl_265});
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2 <= MUX1HOT_s_1_7_2((z_out_1[5]),
          attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_5, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_5,
          apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_5, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_5,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_52_nl, (drf_output_sdt_3_sva_15_0_mx0w3[5]),
          {and_dcpl_257 , operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse ,
          and_dcpl_240 , attention_2_1_16_16_4_4_k_proj_re_or_17_cse , and_dcpl_207
          , and_dcpl_583 , and_dcpl_265});
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3 <= MUX1HOT_s_1_7_2((z_out_1[4]),
          attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_4, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_4,
          apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_4, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_4,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_53_nl, (drf_output_sdt_3_sva_15_0_mx0w3[4]),
          {and_dcpl_257 , operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse ,
          and_dcpl_240 , attention_2_1_16_16_4_4_k_proj_re_or_17_cse , and_dcpl_207
          , and_dcpl_583 , and_dcpl_265});
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4 <= MUX1HOT_s_1_7_2((z_out_1[3]),
          attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_3, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_3,
          apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_3, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_3,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_54_nl, (drf_output_sdt_3_sva_15_0_mx0w3[3]),
          {and_dcpl_257 , operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse ,
          and_dcpl_240 , attention_2_1_16_16_4_4_k_proj_re_or_17_cse , and_dcpl_207
          , and_dcpl_583 , and_dcpl_265});
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5 <= MUX1HOT_s_1_7_2((z_out_1[2]),
          attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_2, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_2,
          apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_2, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_2,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_55_nl, (drf_output_sdt_3_sva_15_0_mx0w3[2]),
          {and_dcpl_257 , operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse ,
          and_dcpl_240 , attention_2_1_16_16_4_4_k_proj_re_or_17_cse , and_dcpl_207
          , and_dcpl_583 , and_dcpl_265});
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6 <= MUX1HOT_s_1_7_2((z_out_1[1]),
          attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_1, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_1,
          apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_1, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_1,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_56_nl, (drf_output_sdt_3_sva_15_0_mx0w3[1]),
          {and_dcpl_257 , operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse ,
          and_dcpl_240 , attention_2_1_16_16_4_4_k_proj_re_or_17_cse , and_dcpl_207
          , and_dcpl_583 , and_dcpl_265});
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7 <= MUX1HOT_s_1_7_2((z_out_1[0]),
          attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_0, RESHAPE_2D_TO_3D_LOOP_3_1_mux_36_cse_0,
          apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_0, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_0_mx0w1_0,
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_57_nl, (drf_output_sdt_3_sva_15_0_mx0w3[0]),
          {and_dcpl_257 , operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_or_3_cse ,
          and_dcpl_240 , attention_2_1_16_16_4_4_k_proj_re_or_17_cse , and_dcpl_207
          , and_dcpl_583 , and_dcpl_265});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_7 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_6 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_5 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_4 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_3 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_2 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_1 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_0 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_15_13 <= 3'b000;
      attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0 <= 13'b0000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_15_8 <= 8'b00000000;
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_7 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_6 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_5 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_4 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_3 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_2 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_1 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_0 <= 1'b0;
      attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_15_0 <= 16'b0000000000000000;
      attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_v_proj_re_and_95_cse ) begin
      attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_0_sva_1_39_16, and_dcpl_1084);
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_1_sva_1_39_16, and_dcpl_1088);
      attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_2_sva_1_39_16, and_dcpl_1091);
      attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_3_sva_1_39_16, and_dcpl_1094);
      attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_4_sva_1_39_16, and_dcpl_1097);
      attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_5_sva_1_39_16, and_dcpl_1100);
      attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_6_sva_1_39_16, and_dcpl_1103);
      attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_7_sva_1_39_16, and_dcpl_1106);
      attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_8_sva_1_39_16, and_dcpl_1109);
      attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_9_sva_1_39_16, and_dcpl_1112);
      attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_10_sva_1_39_16, and_dcpl_1115);
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_11_sva_1_39_16, and_dcpl_1118);
      attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_12_sva_1_39_16, and_dcpl_1121);
      attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_13_sva_1_39_16, and_dcpl_1124);
      attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_14_sva_1_39_16, and_dcpl_1127);
      attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_39_16 <= MUX_v_24_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
          attention_2_1_16_16_4_4_v_proj_re_0_15_sva_1_39_16, and_dcpl_1130);
      attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0, and_dcpl_1084);
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_15_8 <= MUX_v_8_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:8]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8, and_dcpl_1088);
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_7 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[7]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7, and_dcpl_1088);
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_6 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[6]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6, and_dcpl_1088);
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_5 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[5]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5, and_dcpl_1088);
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_4 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[4]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4, and_dcpl_1088);
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_3 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[3]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3, and_dcpl_1088);
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_2 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[2]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2, and_dcpl_1088);
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_1 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[1]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1, and_dcpl_1088);
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_0 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[0]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0, and_dcpl_1088);
      attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_3_0_0_lpi_3_15_0, and_dcpl_1091);
      attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0, and_dcpl_1094);
      attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_3_0_1_lpi_3_15_0, and_dcpl_1097);
      attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_3_0_2_lpi_3_15_0, and_dcpl_1100);
      attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_3_0_3_lpi_3_15_0, and_dcpl_1103);
      attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0, and_dcpl_1106);
      attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_v_proj_re_0_8_lpi_4_15_0, and_dcpl_1109);
      attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_v_proj_re_0_9_lpi_4_15_0, and_dcpl_1112);
      attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_15_13 <= MUX_v_3_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:13]),
          reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd, and_dcpl_1115);
      attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0 <= MUX_v_13_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[12:0]),
          reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1, and_dcpl_1115);
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_15_8 <= MUX_v_8_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:8]),
          apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_15_8, and_dcpl_1118);
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_7 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[7]),
          apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_7, and_dcpl_1118);
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_6 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[6]),
          apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_6, and_dcpl_1118);
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_5 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[5]),
          apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_5, and_dcpl_1118);
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_4 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[4]),
          apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_4, and_dcpl_1118);
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_3 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[3]),
          apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_3, and_dcpl_1118);
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_2 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[2]),
          apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_2, and_dcpl_1118);
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_1 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[1]),
          apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_1, and_dcpl_1118);
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_0 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[0]),
          apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_0, and_dcpl_1118);
      attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0, and_dcpl_1121);
      attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_2_0_1_lpi_3_15_0, and_dcpl_1124);
      attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_2_0_2_lpi_3_15_0, and_dcpl_1127);
      attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0, and_dcpl_1130);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_39_16 <= 24'b000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~(or_dcpl_1146
        | and_dcpl_1055)) ) begin
      attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_39_16 <= attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_39_16 <= 24'b000000000000000000000000;
      attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_15_0 <= 16'b0000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_v_proj_and_30_cse ) begin
      attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_39_16 <= attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16_mx0w5;
      attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_15_0 <= attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0_mx0w6;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva <= 1'b0;
      GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva <= 1'b0;
    end
    else if ( GEMM_3D_FLOAT_LOOP_3_1_and_44_cse ) begin
      GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva <= MUX1HOT_s_1_4_2(APPLY_ROTARY_POS_EMB_LOOP_3_and_7_nl,
          GEMM_3D_FLOAT_LOOP_3_and_tmp_6_sva_mx0w1, GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva_mx0w3,
          (~ QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1),
          {and_dcpl_207 , and_dcpl_1152 , and_dcpl_222 , and_dcpl_1154});
      GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva <= MUX1HOT_s_1_4_2(APPLY_ROTARY_POS_EMB_LOOP_3_and_5_nl,
          GEMM_3D_FLOAT_LOOP_3_and_tmp_7_sva_mx0w1, GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva_mx0w3,
          QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1, {and_dcpl_207
          , and_dcpl_1152 , and_dcpl_222 , and_dcpl_1154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_embed_3_0_3_lpi_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_3_0_2_lpi_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_3_0_1_lpi_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_3_0_0_lpi_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_q_embed_2_0_3_lpi_3 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_q_embed_and_cse ) begin
      attention_2_1_16_16_4_4_q_embed_3_0_3_lpi_3 <= attention_2_1_16_16_4_4_q_embed_mux_14_cse;
      attention_2_1_16_16_4_4_q_embed_3_0_2_lpi_3 <= attention_2_1_16_16_4_4_q_embed_mux_13_cse;
      attention_2_1_16_16_4_4_q_embed_3_0_1_lpi_3 <= attention_2_1_16_16_4_4_q_embed_mux_11_cse;
      attention_2_1_16_16_4_4_q_embed_3_0_0_lpi_3 <= attention_2_1_16_16_4_4_q_embed_mux_9_cse;
      attention_2_1_16_16_4_4_q_embed_2_0_3_lpi_3 <= attention_2_1_16_16_4_4_q_embed_mux_7_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_q_embed_0_0_0_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~((~ mux_2130_nl)
        & and_dcpl_718)) ) begin
      attention_2_1_16_16_4_4_q_embed_0_0_0_sva_1 <= MUX_v_40_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
          attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1, or_dcpl_1025);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_k_embed_0_0_0_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~(mux_2131_nl
        & (~ (fsm_output[8])) & and_dcpl_1145)) ) begin
      attention_2_1_16_16_4_4_k_embed_0_0_0_sva_1 <= apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2_mx0w3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_991)
        | and_dcpl_346 | attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c1
        | and_dcpl_204 | and_dcpl_348 | and_dcpl_349 | and_dcpl_351 | and_dcpl_1162
        | mux_tmp_2153 | attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c9)
        ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          attention_2_1_16_16_4_4_q_embed_mux1h_40_nl, not_4510_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~(or_dcpl_996
        | mux_2159_nl)) | and_dcpl_346 | and_dcpl_204 | and_dcpl_348 | and_dcpl_351
        | mux_tmp_2176 | attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx0c7)
        ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          attention_2_1_16_16_4_4_q_embed_mux1h_41_nl, not_4483_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~(or_dcpl_993
        | mux_2182_nl)) | and_dcpl_346 | and_dcpl_204 | and_dcpl_348 | and_dcpl_351
        | mux_tmp_2176 | attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx0c7)
        ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          attention_2_1_16_16_4_4_q_embed_mux1h_42_nl, not_4482_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_990)
        | and_dcpl_346 | attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c1 |
        and_dcpl_204 | and_dcpl_348 | and_dcpl_349 | and_dcpl_351 | and_dcpl_1162
        | mux_tmp_2153 | attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c9)
        ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          attention_2_1_16_16_4_4_q_embed_mux1h_43_nl, not_4511_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_988)
        | and_dcpl_346 | mux_2198_nl | and_dcpl_204 | and_dcpl_348 | and_dcpl_351
        | mux_tmp_2176 | attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx0c7)
        & (and_dcpl_346 | and_dcpl_204 | and_dcpl_348 | and_dcpl_351 | mux_tmp_2176
        | and_dcpl_352 | attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx0c7)
        ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          attention_2_1_16_16_4_4_q_embed_mux1h_44_nl, not_4512_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_985)
        | and_dcpl_346 | mux_2204_nl | and_dcpl_204 | and_dcpl_348 | and_dcpl_351
        | mux_tmp_2176 | attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx0c7)
        & (and_dcpl_346 | and_dcpl_204 | and_dcpl_348 | and_dcpl_351 | mux_tmp_2176
        | and_dcpl_352 | attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx0c7)
        ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          attention_2_1_16_16_4_4_q_embed_mux1h_45_nl, not_4513_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_980)
        | and_dcpl_346 | mux_2210_nl | and_dcpl_204 | and_dcpl_348 | and_dcpl_351
        | mux_tmp_2176 | attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx0c7)
        & (and_dcpl_346 | and_dcpl_204 | and_dcpl_348 | and_dcpl_351 | mux_tmp_2176
        | and_dcpl_352 | attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx0c7)
        ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          attention_2_1_16_16_4_4_q_embed_mux1h_46_nl, not_4514_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_983)
        | and_dcpl_346 | attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c1 |
        and_dcpl_204 | and_dcpl_348 | and_dcpl_349 | and_dcpl_351 | and_dcpl_1162
        | mux_tmp_2153 | attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c9)
        ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          attention_2_1_16_16_4_4_q_embed_mux1h_47_nl, not_4515_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & ((~ or_dcpl_987)
        | and_dcpl_346 | mux_2226_nl | and_dcpl_204 | and_dcpl_348 | and_dcpl_351
        | mux_tmp_2176 | attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx0c7)
        & (and_dcpl_346 | and_dcpl_204 | and_dcpl_348 | and_dcpl_351 | mux_tmp_2176
        | and_dcpl_352 | attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx0c7)
        ) begin
      attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1 <= MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
          attention_2_1_16_16_4_4_q_embed_mux1h_48_nl, not_4516_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      TRANSPOSE_LAST_TWO_DIMS_LOOP_3_k_2_0_sva_1 <= 3'b000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~((~ (fsm_output[0]))
        | (~ (fsm_output[1])) | (fsm_output[2]) | (~ (fsm_output[4])) | (fsm_output[8])
        | or_dcpl_1134 | (fsm_output[7:6]!=2'b10))) ) begin
      TRANSPOSE_LAST_TWO_DIMS_LOOP_3_k_2_0_sva_1 <= z_out_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_1 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_attn_weights_and_cse ) begin
      attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_35_nl,
          attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2_mx1, and_dcpl_193);
      attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_34_nl,
          attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_2_mx1, and_dcpl_193);
      attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_33_nl,
          attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2_mx1, and_dcpl_193);
      attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_32_nl,
          attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2_mx1, and_dcpl_193);
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_31_nl,
          attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2_mx1, and_dcpl_193);
      attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_30_nl,
          attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2_mx1, and_dcpl_193);
      attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_29_nl,
          attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2_mx1, and_dcpl_193);
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_28_nl,
          attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2_mx1, and_dcpl_193);
      attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_27_nl,
          attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2_mx1, and_dcpl_193);
      attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_26_nl,
          attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2_mx1, and_dcpl_193);
      attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_25_nl,
          attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2_mx1, and_dcpl_193);
      attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_1 <= MUX_v_40_2_2(GEMM_3D_FLOAT_LOOP_3_and_24_nl,
          attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2_mx1, and_dcpl_193);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      GEMM_3D_FLOAT_LOOP_3_and_tmp_sva <= 1'b0;
      GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva <= 1'b0;
      GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva <= 1'b0;
      GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva <= 1'b0;
      GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva <= 1'b0;
      GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva <= 1'b0;
      GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva <= 1'b0;
      GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva <= 1'b0;
    end
    else if ( GEMM_3D_FLOAT_LOOP_3_and_36_cse ) begin
      GEMM_3D_FLOAT_LOOP_3_and_tmp_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_sva_mx0w0;
      GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva_mx0w0;
      GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva_mx0w0;
      GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva_mx0w0;
      GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva_mx0w0;
      GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva_mx0w0;
      GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva_mx0w0;
      GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva <= GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_3 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_attn_weights_and_52_cse ) begin
      attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_6_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1, and_dcpl_1199);
      attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_6_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1, and_dcpl_1199);
      attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_6_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1, and_dcpl_1199);
      attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_6_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1, and_dcpl_1199);
      attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_6_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1, and_dcpl_1199);
      attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_6_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1, and_dcpl_1199);
      attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_6_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1, and_dcpl_1199);
      attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_6_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1, and_dcpl_1199);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_3 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_3 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_attn_weights_and_48_cse ) begin
      attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_6_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx1, and_dcpl_349);
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_6_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx1, and_dcpl_349);
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_6_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx1, and_dcpl_349);
      attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_3 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_6_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx1, and_dcpl_349);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_attn_weights_and_12_cse ) begin
      attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_3,
          attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8_mx1, and_dcpl_377);
      attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1,
          attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9_mx1, and_dcpl_377);
      attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_3,
          attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8_mx1, and_dcpl_377);
      attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_3,
          attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8_mx1, and_dcpl_377);
      attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1,
          attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9_mx1, and_dcpl_377);
      attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_3,
          attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8_mx1, and_dcpl_377);
      attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_3,
          attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8_mx1, and_dcpl_377);
      attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1,
          attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9_mx1, and_dcpl_377);
      attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_3,
          attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8_mx1, and_dcpl_377);
      attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_3,
          attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8_mx1, and_dcpl_377);
      attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1,
          attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9_mx1, and_dcpl_377);
      attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_3,
          attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8_mx1, and_dcpl_377);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_4 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_5 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_4 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_4 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_5 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_4 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_4 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_5 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_4 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_4 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_5 <= 40'b0000000000000000000000000000000000000000;
      attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_4 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_attn_weights_and_24_cse ) begin
      attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx2, and_dcpl_351);
      attention_2_1_16_16_4_4_attn_weights_0_0_0_sva_5 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1_mx2, and_dcpl_351);
      attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx1, and_dcpl_351);
      attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx2, and_dcpl_351);
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_5 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx1, and_dcpl_351);
      attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx2, and_dcpl_351);
      attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx1, and_dcpl_351);
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_5 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx2, and_dcpl_351);
      attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx1, and_dcpl_351);
      attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx1, and_dcpl_351);
      attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_5 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx1, and_dcpl_351);
      attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_4 <= MUX_v_40_2_2(attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8_mx1,
          attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx1, and_dcpl_351);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      softmax_1_4_3_sum_sva_1 <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~(mux_2248_nl
        & and_dcpl_295)) ) begin
      softmax_1_4_3_sum_sva_1 <= softmax_1_4_3_sum_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva <= 1'b0;
      GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva <= 1'b0;
      GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva <= 1'b0;
      GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva <= 1'b0;
    end
    else if ( GEMM_3D_FLOAT_LOOP_3_1_and_46_cse ) begin
      GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva <= GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva_mx0w0;
      GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva <= GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva_mx0w0;
      GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva <= GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva_mx0w0;
      GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva <= GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_abs_4_qr_35_0_lpi_1_dfm_35 <= 1'b0;
      attention_abs_4_qr_35_0_lpi_1_dfm_34_0 <= 35'b00000000000000000000000000000000000;
    end
    else if ( attention_abs_4_qelse_and_ssc ) begin
      attention_abs_4_qr_35_0_lpi_1_dfm_35 <= (attention_abs_qr_35_0_lpi_1_dfm_mx0w0[35])
          & (~ attention_abs_4_qr_35_0_lpi_1_dfm_mx0c1);
      attention_abs_4_qr_35_0_lpi_1_dfm_34_0 <= MUX_v_35_2_2((attention_abs_qr_35_0_lpi_1_dfm_mx0w0[34:0]),
          (operator_40_24_true_AC_TRN_AC_WRAP_operator_40_24_true_AC_TRN_AC_WRAP_acc_psp_sva_1[34:0]),
          attention_abs_4_qr_35_0_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      compute_sqrt_1_guess_sva_34 <= 1'b0;
      compute_sqrt_1_guess_sva_33_0 <= 34'b0000000000000000000000000000000000;
    end
    else if ( compute_sqrt_1_guess_and_ssc ) begin
      compute_sqrt_1_guess_sva_34 <= MUX_s_1_2_2(attention_abs_qr_35_0_lpi_1_dfm_mx1_35,
          (compute_sqrt_1_for_acc_1_itm_40_1_1[34]), and_dcpl_292);
      compute_sqrt_1_guess_sva_33_0 <= MUX_v_34_2_2(attention_abs_qr_35_0_lpi_1_dfm_mx1_34_1,
          (compute_sqrt_1_for_acc_1_itm_40_1_1[33:0]), and_dcpl_292);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_38_0 <= 39'b000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & and_dcpl_548 )
        begin
      QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_38_0 <= QUANTIZE_ACTIVATION_LOOP_1_1_max_val_lpi_2_dfm_1_38_0_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_cse ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
      attention_2_1_16_16_4_4_quantized_final_output_0_1_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_8_cse ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
      attention_2_1_16_16_4_4_quantized_final_output_0_10_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_16_cse ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
      attention_2_1_16_16_4_4_quantized_final_output_0_11_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_24_cse ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
      attention_2_1_16_16_4_4_quantized_final_output_0_12_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_32_cse ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
      attention_2_1_16_16_4_4_quantized_final_output_0_13_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_40_cse ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
      attention_2_1_16_16_4_4_quantized_final_output_0_14_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_48_cse ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
      attention_2_1_16_16_4_4_quantized_final_output_0_2_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_56_cse ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
      attention_2_1_16_16_4_4_quantized_final_output_0_3_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_64_cse ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
      attention_2_1_16_16_4_4_quantized_final_output_0_4_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_72_cse ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
      attention_2_1_16_16_4_4_quantized_final_output_0_5_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_80_cse ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
      attention_2_1_16_16_4_4_quantized_final_output_0_6_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_88_cse ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
      attention_2_1_16_16_4_4_quantized_final_output_0_7_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_96_cse ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
      attention_2_1_16_16_4_4_quantized_final_output_0_8_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_7 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_104_cse ) begin
      reg_attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_0_cse <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_cse;
      attention_2_1_16_16_4_4_quantized_final_output_0_9_sva_1_7 <= RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_and_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~(or_tmp_833 |
        (fsm_output[1:0]!=2'b10) | or_dcpl_1109 | nand_253_cse)) ) begin
      RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva <= z_out_13_71_28[43:4];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~ and_dcpl_414)
        ) begin
      QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva <= LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_7 <= 1'b0;
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3 <= 1'b0;
    end
    else if ( attention_2_1_16_16_4_4_quantized_final_output_and_112_cse ) begin
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_7 <= ~((~ QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1)
          | QUANTIZE_ACTIVATION_LOOP_3_1_nand_seb_1);
      attention_2_1_16_16_4_4_quantized_final_output_0_15_sva_3 <= ~(QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1
          | QUANTIZE_ACTIVATION_LOOP_3_1_nand_seb_1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_0_15_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_0_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_14_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_1_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_13_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_2_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_12_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_3_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_11_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_4_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_10_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_5_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_9_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_6_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_8_sva_1_39_16 <= 24'b000000000000000000000000;
      output_0_7_sva_1_39_16 <= 24'b000000000000000000000000;
    end
    else if ( output_and_16_cse ) begin
      output_0_15_sva_1_39_16 <= output_0_15_lpi_4_39_16_mx1;
      output_0_0_sva_1_39_16 <= output_0_0_lpi_4_39_16_mx1;
      output_0_14_sva_1_39_16 <= output_0_14_lpi_4_39_16_mx1;
      output_0_1_sva_1_39_16 <= output_0_1_lpi_4_39_16_mx1;
      output_0_13_sva_1_39_16 <= output_0_13_lpi_4_39_16_mx1;
      output_0_2_sva_1_39_16 <= output_0_2_lpi_4_39_16_mx1;
      output_0_12_sva_1_39_16 <= output_0_12_lpi_4_39_16_mx1;
      output_0_3_sva_1_39_16 <= output_0_3_lpi_4_39_16_mx1;
      output_0_11_sva_1_39_16 <= output_0_11_lpi_4_39_16_mx1;
      output_0_4_sva_1_39_16 <= output_0_4_lpi_4_39_16_mx1;
      output_0_10_sva_1_39_16 <= output_0_10_lpi_4_39_16_mx1;
      output_0_5_sva_1_39_16 <= output_0_5_lpi_4_39_16_mx1;
      output_0_9_sva_1_39_16 <= output_0_9_lpi_4_39_16_mx1;
      output_0_6_sva_1_39_16 <= output_0_6_lpi_4_39_16_mx1;
      output_0_8_sva_1_39_16 <= output_0_8_lpi_4_39_16_mx1;
      output_0_7_sva_1_39_16 <= output_0_7_lpi_4_39_16_mx1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_mul_mut <= 60'b000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( attention_2_1_16_16_4_4_k_cache_upd_rsc_clken_d_1 & (~(or_dcpl_961
        | or_dcpl_1134 | or_1984_cse)) ) begin
      LINEAR_FORWARD_NO_MUL_LOOP_2_3_mul_mut <= z_out_9;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_0_0_sva_2_29_16 <= 14'b00000000000000;
      output_0_1_sva_2_29_16 <= 14'b00000000000000;
      output_0_2_sva_2_29_16 <= 14'b00000000000000;
      output_0_3_sva_2_29_16 <= 14'b00000000000000;
      output_0_4_sva_2_29_16 <= 14'b00000000000000;
      output_0_5_sva_2_29_16 <= 14'b00000000000000;
      output_0_6_sva_2_29_16 <= 14'b00000000000000;
      output_0_7_sva_2_29_16 <= 14'b00000000000000;
      output_0_8_sva_2_29_16 <= 14'b00000000000000;
      output_0_9_sva_2_29_16 <= 14'b00000000000000;
      output_0_10_sva_2_29_16 <= 14'b00000000000000;
      output_0_11_sva_2_29_16 <= 14'b00000000000000;
      output_0_12_sva_2_29_16 <= 14'b00000000000000;
      output_0_13_sva_2_29_16 <= 14'b00000000000000;
      output_0_14_sva_2_29_16 <= 14'b00000000000000;
      output_0_15_sva_2_29_16 <= 14'b00000000000000;
      output_0_0_sva_2_15_0 <= 16'b0000000000000000;
      output_0_1_sva_2_15_8 <= 8'b00000000;
      output_0_1_sva_2_7 <= 1'b0;
      output_0_1_sva_2_6 <= 1'b0;
      output_0_1_sva_2_5 <= 1'b0;
      output_0_1_sva_2_4 <= 1'b0;
      output_0_1_sva_2_3 <= 1'b0;
      output_0_1_sva_2_2 <= 1'b0;
      output_0_1_sva_2_1 <= 1'b0;
      output_0_1_sva_2_0 <= 1'b0;
      output_0_2_sva_2_15_0 <= 16'b0000000000000000;
      output_0_3_sva_2_15_0 <= 16'b0000000000000000;
      output_0_4_sva_2_15_0 <= 16'b0000000000000000;
      output_0_5_sva_2_15_0 <= 16'b0000000000000000;
      output_0_6_sva_2_15_0 <= 16'b0000000000000000;
      output_0_7_sva_2_15_0 <= 16'b0000000000000000;
      output_0_8_sva_2_15_0 <= 16'b0000000000000000;
      output_0_9_sva_2_15_0 <= 16'b0000000000000000;
      output_0_10_sva_2_15_0 <= 16'b0000000000000000;
      output_0_11_sva_2_15_0 <= 16'b0000000000000000;
      output_0_12_sva_2_15_0 <= 16'b0000000000000000;
      output_0_13_sva_2_15_0 <= 16'b0000000000000000;
      output_0_14_sva_2_15_0 <= 16'b0000000000000000;
      output_0_15_sva_2_15_0 <= 16'b0000000000000000;
    end
    else if ( output_and_64_cse ) begin
      output_0_0_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_0_sva_1_39_16[13:0]), output_and_35_nl);
      output_0_1_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_1_sva_1_39_16[13:0]), output_and_39_nl);
      output_0_2_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_2_sva_1_39_16[13:0]), output_and_43_nl);
      output_0_3_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_3_sva_1_39_16[13:0]), output_and_47_nl);
      output_0_4_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_4_sva_1_39_16[13:0]), output_and_51_nl);
      output_0_5_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_5_sva_1_39_16[13:0]), output_and_55_nl);
      output_0_6_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_6_sva_1_39_16[13:0]), output_and_59_nl);
      output_0_7_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_7_sva_1_39_16[13:0]), output_and_63_nl);
      output_0_8_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_8_sva_1_39_16[13:0]), output_and_61_nl);
      output_0_9_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_9_sva_1_39_16[13:0]), output_and_57_nl);
      output_0_10_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_10_sva_1_39_16[13:0]), output_and_53_nl);
      output_0_11_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_11_sva_1_39_16[13:0]), output_and_49_nl);
      output_0_12_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_12_sva_1_39_16[13:0]), output_and_45_nl);
      output_0_13_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_13_sva_1_39_16[13:0]), output_and_41_nl);
      output_0_14_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_14_sva_1_39_16[13:0]), output_and_37_nl);
      output_0_15_sva_2_29_16 <= MUX_v_14_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[29:16]),
          (output_0_15_sva_1_39_16[13:0]), output_and_33_nl);
      output_0_0_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0, or_dcpl_1155);
      output_0_1_sva_2_15_8 <= MUX_v_8_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:8]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8, or_dcpl_1158);
      output_0_1_sva_2_7 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[7]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7, or_dcpl_1158);
      output_0_1_sva_2_6 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[6]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6, or_dcpl_1158);
      output_0_1_sva_2_5 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[5]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5, or_dcpl_1158);
      output_0_1_sva_2_4 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[4]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4, or_dcpl_1158);
      output_0_1_sva_2_3 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[3]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3, or_dcpl_1158);
      output_0_1_sva_2_2 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[2]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2, or_dcpl_1158);
      output_0_1_sva_2_1 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[1]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1, or_dcpl_1158);
      output_0_1_sva_2_0 <= MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[0]),
          APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0, or_dcpl_1158);
      output_0_2_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0, or_dcpl_1160);
      output_0_3_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0, or_dcpl_1162);
      output_0_4_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0, or_dcpl_1165);
      output_0_5_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0, or_dcpl_1167);
      output_0_6_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0, or_dcpl_1169);
      output_0_7_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0, or_dcpl_1141);
      output_0_8_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0, or_dcpl_1170);
      output_0_9_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0, or_dcpl_1168);
      output_0_10_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0, or_dcpl_1166);
      output_0_11_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0, or_dcpl_1164);
      output_0_12_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0, or_dcpl_1161);
      output_0_13_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0, or_dcpl_1159);
      output_0_14_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0, or_dcpl_1156);
      output_0_15_sva_2_15_0 <= MUX_v_16_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
          attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0, or_dcpl_1152);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd <= 1'b0;
      reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 <= 1'b0;
    end
    else if ( GEMM_3D_FLOAT_LOOP_4_l_and_ssc ) begin
      reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd <= GEMM_3D_FLOAT_LOOP_4_l_mux1h_6_nl
          & (~ GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c2);
      reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 <= GEMM_3D_FLOAT_LOOP_4_l_mux1h_8_nl
          & (~ GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c2);
    end
  end
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_nl = MUX1HOT_v_8_4_2((drf_output_sdt_2_sva_15_0_mx0w0[15:8]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd, (drf_output_sdt_3_sva_15_0_mx0w3[15:8]),
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_265 , and_dcpl_268});
  assign not_4947_nl = ~ or_dcpl_1048;
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_1_nl = MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0[7]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7, (drf_output_sdt_3_sva_15_0_mx0w3[7]),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_265 , and_dcpl_268});
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_2_nl = MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0[6]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6, (drf_output_sdt_3_sva_15_0_mx0w3[6]),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_265 , and_dcpl_268});
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_3_nl = MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0[5]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5, (drf_output_sdt_3_sva_15_0_mx0w3[5]),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_265 , and_dcpl_268});
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_4_nl = MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0[4]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4, (drf_output_sdt_3_sva_15_0_mx0w3[4]),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_265 , and_dcpl_268});
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_5_nl = MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0[3]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3, (drf_output_sdt_3_sva_15_0_mx0w3[3]),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_265 , and_dcpl_268});
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_6_nl = MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0[2]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2, (drf_output_sdt_3_sva_15_0_mx0w3[2]),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_265 , and_dcpl_268});
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_7_nl = MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0[1]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1, (drf_output_sdt_3_sva_15_0_mx0w3[1]),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_265 , and_dcpl_268});
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_2_mux1h_8_nl = MUX1HOT_s_1_4_2((drf_output_sdt_2_sva_15_0_mx0w0[0]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0, (drf_output_sdt_3_sva_15_0_mx0w3[0]),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_265 , and_dcpl_268});
  assign rms_norm_16_mux1h_nl = MUX1HOT_s_1_5_2(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4,
      (compute_sqrt_for_acc_1_itm_40_1_1[39]), attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_39,
      reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd, (compute_sqrt_1_for_acc_1_itm_40_1_1[39]),
      {and_321_ssc , and_dcpl_290 , and_dcpl_276 , and_dcpl_278 , and_dcpl_292});
  assign rms_norm_16_mux1h_9_nl = MUX1HOT_v_4_5_2(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0,
      (compute_sqrt_for_acc_1_itm_40_1_1[38:35]), (attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_38_0[38:35]),
      (reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[38:35]), (compute_sqrt_1_for_acc_1_itm_40_1_1[38:35]),
      {and_321_ssc , and_dcpl_290 , and_dcpl_276 , and_dcpl_278 , and_dcpl_292});
  assign operator_40_24_true_AC_TRN_AC_WRAP_1_not_1_nl = ~ mux_851_ssc;
  assign SOFTMAX_LOOP_5_mux_24_nl = MUX_s_1_2_2((SOFTMAX_LOOP_5_mux_12_psp_mx0w0[39]),
      reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd, and_329_ssc);
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_2_mux1h_2_nl = MUX1HOT_v_24_4_2(LINEAR_FORWARD_NO_MUL_LOOP_2_2_conc_1_mut_71_48_mx0w0,
      for_for_strm_in_tmp_sva_25_2, LINEAR_FORWARD_NO_MUL_LOOP_2_3_conc_1_mut_71_48_mx0w3,
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_265 , and_dcpl_268});
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_2_not_nl = ~ or_dcpl_1048;
  assign mux_862_nl = MUX_s_1_2_2((~ mux_tmp_787), or_1732_cse, for_for_and_tmp);
  assign rms_norm_16_mux1h_10_nl = MUX1HOT_s_1_4_2((compute_sqrt_for_acc_1_itm_40_1_1[0]),
      (reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[0]), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut_mx0w2[0]),
      (LINEAR_FORWARD_NO_MUL_LOOP_2_1_mul_mut[0]), {and_dcpl_290 , and_343_itm ,
      and_dcpl_257 , and_dcpl_260});
  assign rms_norm_16_mux1h_6_nl = MUX1HOT_v_24_3_2(LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48_mx0w2,
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48, APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16,
      {and_dcpl_257 , and_dcpl_260 , and_dcpl_310});
  assign rms_norm_16_not_nl = ~ rms_norm_16_div_cmp_a_mx0c0;
  assign rms_norm_16_mux1h_7_nl = MUX1HOT_v_8_3_2((z_out_1[15:8]), LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_310});
  assign rms_norm_16_not_1_nl = ~ rms_norm_16_div_cmp_a_mx0c0;
  assign rms_norm_16_mux1h_11_nl = MUX1HOT_s_1_3_2((z_out_1[7]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_310});
  assign rms_norm_16_mux1h_13_nl = MUX1HOT_s_1_3_2((z_out_1[6]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_310});
  assign rms_norm_16_mux1h_14_nl = MUX1HOT_s_1_3_2((z_out_1[5]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_310});
  assign rms_norm_16_mux1h_15_nl = MUX1HOT_s_1_3_2((z_out_1[4]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_310});
  assign rms_norm_16_mux1h_16_nl = MUX1HOT_s_1_3_2((z_out_1[3]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_310});
  assign rms_norm_16_mux1h_17_nl = MUX1HOT_s_1_3_2((z_out_1[2]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_310});
  assign rms_norm_16_mux1h_18_nl = MUX1HOT_s_1_3_2((z_out_1[1]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_310});
  assign rms_norm_16_mux1h_19_nl = MUX1HOT_s_1_3_2((z_out_1[0]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0, {and_dcpl_257 , and_dcpl_260
      , and_dcpl_310});
  assign INIT_2D_MEM_LOOP_2_mux_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_633_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_nl = INIT_2D_MEM_LOOP_2_mux_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_10_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_6,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_633_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_38_nl = INIT_2D_MEM_LOOP_2_mux_10_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_11_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_5,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_633_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_39_nl = INIT_2D_MEM_LOOP_2_mux_11_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_12_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_4,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_633_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_40_nl = INIT_2D_MEM_LOOP_2_mux_12_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_13_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_3,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_633_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_41_nl = INIT_2D_MEM_LOOP_2_mux_13_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_14_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_2,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_633_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_42_nl = INIT_2D_MEM_LOOP_2_mux_14_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_15_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_1,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_633_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_43_nl = INIT_2D_MEM_LOOP_2_mux_15_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_16_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_1_lpi_3_0,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_633_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_44_nl = INIT_2D_MEM_LOOP_2_mux_16_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_1_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_654_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_1_nl = INIT_2D_MEM_LOOP_2_mux_1_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_17_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_6,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_654_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_24_nl = INIT_2D_MEM_LOOP_2_mux_17_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_18_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_5,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_654_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_25_nl = INIT_2D_MEM_LOOP_2_mux_18_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_19_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_4,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_654_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_26_nl = INIT_2D_MEM_LOOP_2_mux_19_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_20_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_3,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_654_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_27_nl = INIT_2D_MEM_LOOP_2_mux_20_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_21_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_2,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_654_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_28_nl = INIT_2D_MEM_LOOP_2_mux_21_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_22_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_1,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_654_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_29_nl = INIT_2D_MEM_LOOP_2_mux_22_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_23_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_2_lpi_3_0,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_654_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_30_nl = INIT_2D_MEM_LOOP_2_mux_23_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_2_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_648_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_2_nl = INIT_2D_MEM_LOOP_2_mux_2_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_24_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_6,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_648_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_10_nl = INIT_2D_MEM_LOOP_2_mux_24_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_25_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_5,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_648_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_11_nl = INIT_2D_MEM_LOOP_2_mux_25_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_26_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_4,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_648_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_12_nl = INIT_2D_MEM_LOOP_2_mux_26_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_27_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_3,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_648_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_13_nl = INIT_2D_MEM_LOOP_2_mux_27_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_28_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_2,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_648_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_14_nl = INIT_2D_MEM_LOOP_2_mux_28_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_29_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_1,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_648_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_15_nl = INIT_2D_MEM_LOOP_2_mux_29_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_30_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_1_0_3_lpi_3_0,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_648_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_16_nl = INIT_2D_MEM_LOOP_2_mux_30_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_3_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_642_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_3_nl = INIT_2D_MEM_LOOP_2_mux_3_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_31_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_6,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_642_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_17_nl = INIT_2D_MEM_LOOP_2_mux_31_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_32_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_5,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_642_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_18_nl = INIT_2D_MEM_LOOP_2_mux_32_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_33_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_4,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_642_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_19_nl = INIT_2D_MEM_LOOP_2_mux_33_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_34_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_3,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_642_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_20_nl = INIT_2D_MEM_LOOP_2_mux_34_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_35_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_2,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_642_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_21_nl = INIT_2D_MEM_LOOP_2_mux_35_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_36_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_1,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_642_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_22_nl = INIT_2D_MEM_LOOP_2_mux_36_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_37_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_0_lpi_3_0,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_642_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_23_nl = INIT_2D_MEM_LOOP_2_mux_37_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_4_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_636_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_4_nl = INIT_2D_MEM_LOOP_2_mux_4_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_38_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_6,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_636_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_31_nl = INIT_2D_MEM_LOOP_2_mux_38_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_39_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_5,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_636_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_32_nl = INIT_2D_MEM_LOOP_2_mux_39_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_40_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_4,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_636_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_33_nl = INIT_2D_MEM_LOOP_2_mux_40_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_41_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_3,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_636_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_34_nl = INIT_2D_MEM_LOOP_2_mux_41_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_42_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_2,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_636_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_35_nl = INIT_2D_MEM_LOOP_2_mux_42_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_43_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_1,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_636_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_36_nl = INIT_2D_MEM_LOOP_2_mux_43_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_44_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_1_lpi_3_0,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_636_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_37_nl = INIT_2D_MEM_LOOP_2_mux_44_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_5_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_629_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_5_nl = INIT_2D_MEM_LOOP_2_mux_5_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_45_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_6,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_629_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_45_nl = INIT_2D_MEM_LOOP_2_mux_45_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_46_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_5,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_629_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_46_nl = INIT_2D_MEM_LOOP_2_mux_46_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_47_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_4,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_629_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_47_nl = INIT_2D_MEM_LOOP_2_mux_47_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_48_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_3,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_629_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_48_nl = INIT_2D_MEM_LOOP_2_mux_48_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_49_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_2,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_629_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_49_nl = INIT_2D_MEM_LOOP_2_mux_49_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_50_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_1,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_629_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_50_nl = INIT_2D_MEM_LOOP_2_mux_50_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_51_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_2_0_2_lpi_3_0,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_629_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_51_nl = INIT_2D_MEM_LOOP_2_mux_51_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_6_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_639_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_6_nl = INIT_2D_MEM_LOOP_2_mux_6_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_52_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_6,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_639_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_52_nl = INIT_2D_MEM_LOOP_2_mux_52_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_53_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_5,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_639_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_53_nl = INIT_2D_MEM_LOOP_2_mux_53_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_54_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_4,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_639_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_54_nl = INIT_2D_MEM_LOOP_2_mux_54_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_55_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_3,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_639_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_55_nl = INIT_2D_MEM_LOOP_2_mux_55_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_56_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_2,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_639_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_56_nl = INIT_2D_MEM_LOOP_2_mux_56_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_57_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_1,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_639_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_57_nl = INIT_2D_MEM_LOOP_2_mux_57_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_58_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_0_lpi_3_0,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_639_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_58_nl = INIT_2D_MEM_LOOP_2_mux_58_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_7_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_645_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_7_nl = INIT_2D_MEM_LOOP_2_mux_7_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_59_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_6,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_645_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_59_nl = INIT_2D_MEM_LOOP_2_mux_59_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_60_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_5,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_645_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_60_nl = INIT_2D_MEM_LOOP_2_mux_60_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_61_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_4,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_645_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_61_nl = INIT_2D_MEM_LOOP_2_mux_61_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_62_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_3,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_645_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_62_nl = INIT_2D_MEM_LOOP_2_mux_62_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_63_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_2,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_645_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_63_nl = INIT_2D_MEM_LOOP_2_mux_63_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_64_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_1,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_645_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_64_nl = INIT_2D_MEM_LOOP_2_mux_64_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_65_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_1_lpi_3_0,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_645_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_65_nl = INIT_2D_MEM_LOOP_2_mux_65_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_8_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_651_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_8_nl = INIT_2D_MEM_LOOP_2_mux_8_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_66_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_6,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_651_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_66_nl = INIT_2D_MEM_LOOP_2_mux_66_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_67_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_5,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_651_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_67_nl = INIT_2D_MEM_LOOP_2_mux_67_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_68_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_4,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_651_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_68_nl = INIT_2D_MEM_LOOP_2_mux_68_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_69_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_3,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_651_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_69_nl = INIT_2D_MEM_LOOP_2_mux_69_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_70_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_2,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_651_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_70_nl = INIT_2D_MEM_LOOP_2_mux_70_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_71_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_1,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_651_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_71_nl = INIT_2D_MEM_LOOP_2_mux_71_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_72_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_2_lpi_3_0,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_651_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_72_nl = INIT_2D_MEM_LOOP_2_mux_72_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_9_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_7,
      QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1, and_657_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_9_nl = INIT_2D_MEM_LOOP_2_mux_9_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_73_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_6,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_657_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_73_nl = INIT_2D_MEM_LOOP_2_mux_73_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_74_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_5,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_657_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_74_nl = INIT_2D_MEM_LOOP_2_mux_74_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_75_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_4,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_657_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_75_nl = INIT_2D_MEM_LOOP_2_mux_75_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_76_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_3,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_657_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_76_nl = INIT_2D_MEM_LOOP_2_mux_76_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_77_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_2,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_657_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_77_nl = INIT_2D_MEM_LOOP_2_mux_77_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_78_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_1,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_657_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_78_nl = INIT_2D_MEM_LOOP_2_mux_78_nl
      & (~ or_dcpl_1104);
  assign INIT_2D_MEM_LOOP_2_mux_79_nl = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_3_0_3_lpi_3_0,
      (~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1), and_657_itm);
  assign INIT_2D_MEM_LOOP_2_INIT_2D_MEM_LOOP_2_and_79_nl = INIT_2D_MEM_LOOP_2_mux_79_nl
      & (~ or_dcpl_1104);
  assign and_779_nl = and_dcpl_732 & and_dcpl_730;
  assign and_1653_nl = (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd) &
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2==2'b11);
  assign mux_1556_nl = MUX_s_1_2_2(mux_1555_cse, mux_1553_cse, and_1653_nl);
  assign mux_1558_nl = MUX_s_1_2_2(mux_1557_cse, mux_1556_nl, fsm_output[0]);
  assign mux_1560_nl = MUX_s_1_2_2(mux_1559_cse, mux_1558_nl, and_1773_cse);
  assign mux_1561_nl = MUX_s_1_2_2(mux_1560_nl, mux_1546_cse, fsm_output[7]);
  assign and_783_nl = and_dcpl_736 & and_dcpl_730;
  assign and_790_nl = and_dcpl_743 & and_dcpl_740 & and_dcpl_728;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_5_nl = MUX1HOT_v_16_5_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0, (rms_norm_16_div_cmp_z_oreg[15:0]),
      output_0_7_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3, {and_779_nl , (~ mux_1561_nl)
      , and_783_nl , and_dcpl_739 , and_790_nl});
  assign not_4472_nl = ~ and_dcpl_619;
  assign and_943_nl = and_dcpl_732 & and_dcpl_842;
  assign nor_466_nl = ~((~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd)
      | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b10));
  assign mux_1655_nl = MUX_s_1_2_2(mux_1555_cse, mux_1553_cse, nor_466_nl);
  assign mux_1657_nl = MUX_s_1_2_2(mux_1557_cse, mux_1655_nl, fsm_output[0]);
  assign mux_1659_nl = MUX_s_1_2_2(mux_1559_cse, mux_1657_nl, and_1773_cse);
  assign mux_1660_nl = MUX_s_1_2_2(mux_1659_nl, mux_1645_cse, fsm_output[7]);
  assign attention_2_1_16_16_4_4_k_proj_re_nand_nl = ~(mux_1660_nl & (~(or_dcpl_1010
      & and_dcpl_207)));
  assign attention_2_1_16_16_4_4_k_proj_re_and_81_nl = (~ or_dcpl_1010) & and_dcpl_207;
  assign and_945_nl = and_dcpl_743 & and_dcpl_551 & and_dcpl_841;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_30_nl = MUX1HOT_v_16_7_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0, (rms_norm_16_div_cmp_z_oreg[15:0]),
      RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_15_0, output_0_10_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      {and_943_nl , attention_2_1_16_16_4_4_k_proj_re_nand_nl , and_dcpl_843 , attention_2_1_16_16_4_4_k_proj_re_and_81_nl
      , and_dcpl_847 , and_dcpl_739 , and_945_nl});
  assign not_4469_nl = ~ and_dcpl_619;
  assign and_946_nl = and_dcpl_732 & and_dcpl_855;
  assign and_1684_nl = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & (~
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1) & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2==2'b11);
  assign mux_1671_nl = MUX_s_1_2_2(mux_1555_cse, mux_1553_cse, and_1684_nl);
  assign mux_1673_nl = MUX_s_1_2_2(mux_1557_cse, mux_1671_nl, fsm_output[0]);
  assign mux_1675_nl = MUX_s_1_2_2(mux_1559_cse, mux_1673_nl, and_1773_cse);
  assign mux_1676_nl = MUX_s_1_2_2(mux_1675_nl, mux_1645_cse, fsm_output[7]);
  assign attention_2_1_16_16_4_4_k_proj_re_nand_2_nl = ~(mux_1676_nl & (~(or_dcpl_1012
      & and_dcpl_207)));
  assign attention_2_1_16_16_4_4_k_proj_re_and_83_nl = (~ or_dcpl_1012) & and_dcpl_207;
  assign and_948_nl = and_dcpl_743 & and_dcpl_551 & and_dcpl_854;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_32_nl = MUX1HOT_v_16_7_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0, (rms_norm_16_div_cmp_z_oreg[15:0]),
      RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_15_0, output_0_11_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      {and_946_nl , attention_2_1_16_16_4_4_k_proj_re_nand_2_nl , and_dcpl_856 ,
      attention_2_1_16_16_4_4_k_proj_re_and_83_nl , and_dcpl_847 , and_dcpl_739 ,
      and_948_nl});
  assign not_4468_nl = ~ and_dcpl_619;
  assign and_949_nl = and_dcpl_732 & and_dcpl_859;
  assign or_2589_nl = (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd) |
      (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1) | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b00);
  assign mux_1687_nl = MUX_s_1_2_2(mux_1553_cse, mux_1555_cse, or_2589_nl);
  assign mux_1689_nl = MUX_s_1_2_2(mux_1557_cse, mux_1687_nl, fsm_output[0]);
  assign mux_1691_nl = MUX_s_1_2_2(mux_1559_cse, mux_1689_nl, and_1773_cse);
  assign mux_1692_nl = MUX_s_1_2_2(mux_1691_nl, mux_1645_cse, fsm_output[7]);
  assign attention_2_1_16_16_4_4_k_proj_re_nand_4_nl = ~(mux_1692_nl & (~(or_dcpl_1014
      & and_dcpl_207)));
  assign attention_2_1_16_16_4_4_k_proj_re_and_85_nl = (~ or_dcpl_1014) & and_dcpl_207;
  assign and_951_nl = and_dcpl_743 & and_dcpl_740 & and_dcpl_818;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_34_nl = MUX1HOT_v_16_7_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0, (rms_norm_16_div_cmp_z_oreg[15:0]),
      RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_15_0, output_0_12_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      {and_949_nl , attention_2_1_16_16_4_4_k_proj_re_nand_4_nl , and_dcpl_860 ,
      attention_2_1_16_16_4_4_k_proj_re_and_85_nl , and_dcpl_847 , and_dcpl_739 ,
      and_951_nl});
  assign not_4467_nl = ~ and_dcpl_619;
  assign and_952_nl = and_dcpl_732 & and_dcpl_863;
  assign nand_367_nl = ~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2==2'b01));
  assign mux_1703_nl = MUX_s_1_2_2(mux_1553_cse, mux_1555_cse, nand_367_nl);
  assign mux_1705_nl = MUX_s_1_2_2(mux_1557_cse, mux_1703_nl, fsm_output[0]);
  assign mux_1707_nl = MUX_s_1_2_2(mux_1559_cse, mux_1705_nl, and_1773_cse);
  assign mux_1708_nl = MUX_s_1_2_2(mux_1707_nl, mux_1645_cse, fsm_output[7]);
  assign attention_2_1_16_16_4_4_k_proj_re_nand_6_nl = ~(mux_1708_nl & (~(or_dcpl_1016
      & and_dcpl_207)));
  assign attention_2_1_16_16_4_4_k_proj_re_and_87_nl = (~ or_dcpl_1016) & and_dcpl_207;
  assign and_954_nl = and_dcpl_743 & and_dcpl_740 & and_dcpl_830;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_36_nl = MUX1HOT_v_16_7_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0, (rms_norm_16_div_cmp_z_oreg[15:0]),
      RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_15_0, output_0_13_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      {and_952_nl , attention_2_1_16_16_4_4_k_proj_re_nand_6_nl , and_dcpl_864 ,
      attention_2_1_16_16_4_4_k_proj_re_and_87_nl , and_dcpl_847 , and_dcpl_739 ,
      and_954_nl});
  assign not_4466_nl = ~ and_dcpl_619;
  assign and_955_nl = and_dcpl_732 & and_dcpl_871;
  assign and_1697_nl = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2==2'b10);
  assign mux_1719_nl = MUX_s_1_2_2(mux_1555_cse, mux_1553_cse, and_1697_nl);
  assign mux_1721_nl = MUX_s_1_2_2(mux_1557_cse, mux_1719_nl, fsm_output[0]);
  assign mux_1723_nl = MUX_s_1_2_2(mux_1559_cse, mux_1721_nl, and_1773_cse);
  assign mux_1724_nl = MUX_s_1_2_2(mux_1723_nl, mux_1645_cse, fsm_output[7]);
  assign attention_2_1_16_16_4_4_k_proj_re_nand_8_nl = ~(mux_1724_nl & (~(or_dcpl_1018
      & and_dcpl_207)));
  assign attention_2_1_16_16_4_4_k_proj_re_and_89_nl = (~ or_dcpl_1018) & and_dcpl_207;
  assign and_957_nl = and_dcpl_743 & and_dcpl_740 & and_dcpl_841;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_38_nl = MUX1HOT_v_16_7_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0, (rms_norm_16_div_cmp_z_oreg[15:0]),
      RESHAPE_2D_TO_3D_LOOP_3_2_slc_attention_2_1_16_16_4_4_v_proj_re_40_39_0_ctmp_sva_15_0_1,
      attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_15_0, output_0_14_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      {and_955_nl , attention_2_1_16_16_4_4_k_proj_re_nand_8_nl , and_dcpl_872 ,
      attention_2_1_16_16_4_4_k_proj_re_and_89_nl , and_dcpl_847 , and_dcpl_739 ,
      and_957_nl});
  assign not_4465_nl = ~ and_dcpl_619;
  assign and_960_nl = and_dcpl_732 & and_dcpl_850;
  assign or_2611_nl = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd | (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1)
      | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b00);
  assign mux_1738_nl = MUX_s_1_2_2(mux_1553_cse, mux_1555_cse, or_2611_nl);
  assign mux_1740_nl = MUX_s_1_2_2(mux_1557_cse, mux_1738_nl, fsm_output[0]);
  assign mux_1742_nl = MUX_s_1_2_2(mux_1559_cse, mux_1740_nl, and_1773_cse);
  assign mux_1743_nl = MUX_s_1_2_2(mux_1742_nl, mux_1546_cse, fsm_output[7]);
  assign and_962_nl = and_dcpl_743 & and_dcpl_740 & and_dcpl_550;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_42_nl = MUX1HOT_v_16_5_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0, (rms_norm_16_div_cmp_z_oreg[15:0]),
      output_0_4_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3, {and_960_nl , (~ mux_1743_nl)
      , and_dcpl_851 , and_dcpl_739 , and_962_nl});
  assign not_4463_nl = ~ and_dcpl_619;
  assign and_963_nl = and_dcpl_732 & and_dcpl_836;
  assign or_2617_nl = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd | (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1)
      | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b01);
  assign mux_1754_nl = MUX_s_1_2_2(mux_1553_cse, mux_1555_cse, or_2617_nl);
  assign mux_1756_nl = MUX_s_1_2_2(mux_1557_cse, mux_1754_nl, fsm_output[0]);
  assign mux_1758_nl = MUX_s_1_2_2(mux_1559_cse, mux_1756_nl, and_1773_cse);
  assign mux_1759_nl = MUX_s_1_2_2(mux_1758_nl, mux_1546_cse, fsm_output[7]);
  assign and_965_nl = and_dcpl_743 & and_dcpl_740 & and_dcpl_835;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_44_nl = MUX1HOT_v_16_5_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0, (rms_norm_16_div_cmp_z_oreg[15:0]),
      output_0_5_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3, {and_963_nl , (~ mux_1759_nl)
      , and_dcpl_837 , and_dcpl_739 , and_965_nl});
  assign not_4462_nl = ~ and_dcpl_619;
  assign and_966_nl = and_dcpl_732 & and_dcpl_826;
  assign nor_500_nl = ~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd | (~
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1) | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b10));
  assign mux_1770_nl = MUX_s_1_2_2(mux_1555_cse, mux_1553_cse, nor_500_nl);
  assign mux_1772_nl = MUX_s_1_2_2(mux_1557_cse, mux_1770_nl, fsm_output[0]);
  assign mux_1774_nl = MUX_s_1_2_2(mux_1559_cse, mux_1772_nl, and_1773_cse);
  assign mux_1775_nl = MUX_s_1_2_2(mux_1774_nl, mux_1546_cse, fsm_output[7]);
  assign and_968_nl = and_dcpl_743 & and_dcpl_740 & and_dcpl_825;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_46_nl = MUX1HOT_v_16_5_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0, (rms_norm_16_div_cmp_z_oreg[15:0]),
      output_0_6_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3, {and_966_nl , (~ mux_1775_nl)
      , and_dcpl_827 , and_dcpl_739 , and_968_nl});
  assign not_4461_nl = ~ and_dcpl_619;
  assign and_969_nl = and_dcpl_732 & and_dcpl_820;
  assign or_2492_nl = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b00)
      | (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd) | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  assign mux_1786_nl = MUX_s_1_2_2(mux_1553_cse, mux_1555_cse, or_2492_nl);
  assign mux_1788_nl = MUX_s_1_2_2(mux_1557_cse, mux_1786_nl, fsm_output[0]);
  assign mux_1790_nl = MUX_s_1_2_2(mux_1559_cse, mux_1788_nl, and_1773_cse);
  assign mux_1791_nl = MUX_s_1_2_2(mux_1790_nl, mux_1546_cse, fsm_output[7]);
  assign and_971_nl = and_dcpl_743 & and_dcpl_551 & and_dcpl_818;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_48_nl = MUX1HOT_v_16_5_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0, (rms_norm_16_div_cmp_z_oreg[15:0]),
      output_0_8_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3, {and_969_nl , (~ mux_1791_nl)
      , and_dcpl_821 , and_dcpl_739 , and_971_nl});
  assign not_4460_nl = ~ and_dcpl_619;
  assign and_972_nl = and_dcpl_732 & and_dcpl_831;
  assign or_2497_nl = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b01)
      | (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd) | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  assign mux_1802_nl = MUX_s_1_2_2(mux_1553_cse, mux_1555_cse, or_2497_nl);
  assign mux_1804_nl = MUX_s_1_2_2(mux_1557_cse, mux_1802_nl, fsm_output[0]);
  assign mux_1806_nl = MUX_s_1_2_2(mux_1559_cse, mux_1804_nl, and_1773_cse);
  assign mux_1807_nl = MUX_s_1_2_2(mux_1806_nl, mux_1546_cse, fsm_output[7]);
  assign and_974_nl = and_dcpl_743 & and_dcpl_551 & and_dcpl_830;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_50_nl = MUX1HOT_v_16_5_2(z_out_1,
      attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0, (rms_norm_16_div_cmp_z_oreg[15:0]),
      output_0_9_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3, {and_972_nl , (~ mux_1807_nl)
      , and_dcpl_832 , and_dcpl_739 , and_974_nl});
  assign not_4459_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_68_nl = MUX1HOT_v_8_6_2((z_out_1[15:8]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0[15:8]), (rms_norm_16_div_cmp_z_oreg[15:8]),
      APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8,
      (output_0_2_lpi_3_15_0[15:8]), (drf_output_sdt_3_sva_15_0_mx0w3[15:8]), {and_1034_itm
      , (~ mux_1966_itm) , and_dcpl_989 , and_dcpl_374 , and_dcpl_739 , and_1037_itm});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_118_nl = MUX1HOT_v_8_6_2((z_out_1[7:0]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0[7:0]), (rms_norm_16_div_cmp_z_oreg[7:0]),
      ({APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7
      , APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6
      , APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5
      , APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4
      , APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3
      , APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2
      , APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1
      , APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0}),
      (output_0_2_lpi_3_15_0[7:0]), (drf_output_sdt_3_sva_15_0_mx0w3[7:0]), {and_1034_itm
      , (~ mux_1966_itm) , and_dcpl_989 , and_dcpl_374 , and_dcpl_739 , and_1037_itm});
  assign not_4443_nl = ~ and_dcpl_619;
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_39_nl = MUX_v_24_16_2(({reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd
      , (reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[38:16])}), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[39:16]),
      apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_39_16, apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16,
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3[39:16]), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm[39:16]),
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_39_16, apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_39_16,
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3[39:16]), (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm[39:16]),
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_39_16, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16,
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3[39:16]), (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm[39:16]),
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_39_16, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_58_nl = MUX1HOT_v_24_7_2(attention_2_1_16_16_4_4_v_proj_re_0_12_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_39_16,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16_mx0w1, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16_mx0w1,
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_39_16, APPLY_ROTARY_POS_EMB_LOOP_6_mux_39_nl,
      {and_dcpl_726 , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207
      , and_dcpl_847 , and_dcpl_583});
  assign not_4582_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_59_nl = MUX1HOT_v_24_6_2(attention_2_1_16_16_4_4_v_proj_re_0_14_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16_mx0w1, apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16_mx0w1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16, {and_dcpl_726
      , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign not_4583_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_60_nl = MUX1HOT_v_24_6_2(attention_2_1_16_16_4_4_v_proj_re_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16_mx0w1, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16_mx0w1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16, {and_dcpl_726
      , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign not_4584_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_61_nl = MUX1HOT_v_24_6_2(attention_2_1_16_16_4_4_v_proj_re_0_5_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_39_16, attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_1_0_3_lpi_3_39_16_mx0w5,
      attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_39_16, {and_dcpl_726 , and_dcpl_983
      , and_dcpl_240 , and_dcpl_626 , and_dcpl_207 , and_dcpl_213});
  assign not_4585_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_62_nl = MUX1HOT_v_24_6_2(attention_2_1_16_16_4_4_v_proj_re_0_6_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_39_16_mx0w1, {and_dcpl_726 , attention_2_1_16_16_4_4_k_proj_re_or_cse
      , and_dcpl_983 , and_dcpl_240 , attention_2_1_16_16_4_4_k_proj_re_or_17_cse
      , and_dcpl_207});
  assign not_4586_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_63_nl = MUX1HOT_v_24_6_2(attention_2_1_16_16_4_4_v_proj_re_0_8_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_39_16, {and_dcpl_726 , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign not_4587_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_64_nl = MUX1HOT_v_24_6_2(attention_2_1_16_16_4_4_v_proj_re_0_9_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16_mx0w1, attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_39_16, {and_dcpl_726 , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign not_4588_nl = ~ and_dcpl_619;
  assign APPLY_ROTARY_POS_EMB_LOOP_3_APPLY_ROTARY_POS_EMB_LOOP_3_nor_nl = ~(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_or_2_nl = and_dcpl_1151
      | compute_sqrt_for_i_and_2_cse;
  assign QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_1_nl = MUX1HOT_s_1_6_2((LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_2[0]),
      APPLY_ROTARY_POS_EMB_LOOP_3_APPLY_ROTARY_POS_EMB_LOOP_3_nor_nl, LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0,
      GEMM_3D_FLOAT_LOOP_3_and_tmp_4_sva_mx0w2, GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_0_sva_mx0w3,
      (~ QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1), {and_dcpl_725
      , RMS_NORM_LOOP_2_2_i_and_9_cse , QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_or_2_nl
      , and_dcpl_1152 , and_dcpl_222 , and_dcpl_557});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_95_nl = MUX_v_2_2_2((reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1[12:11]),
      2'b10, and_dcpl_1363);
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_96_nl = MUX_s_1_2_2((reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1[10]),
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1, and_dcpl_1363);
  assign APPLY_ROTARY_POS_EMB_LOOP_6_APPLY_ROTARY_POS_EMB_LOOP_6_or_7_nl = (reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1[9])
      | and_dcpl_1363;
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_97_nl = MUX_s_1_2_2((reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1[8]),
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2,
      and_dcpl_1363);
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_98_nl = MUX_v_8_2_2((reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1[7:0]),
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3,
      and_dcpl_1363);
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_99_nl = MUX_v_24_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_39_16,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[39:16]), and_dcpl_1363);
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_100_nl = MUX_v_8_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[15:8]), and_dcpl_1363);
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_101_nl = MUX_v_8_2_2(({APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6 , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4 , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2 , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0}), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[7:0]),
      and_dcpl_1363);
  assign nl_APPLY_ROTARY_POS_EMB_LOOP_6_mul_3_itm  = $signed(conv_u2s_16_17(signext_16_14({(~
      and_dcpl_1363) , APPLY_ROTARY_POS_EMB_LOOP_6_mux_95_nl , APPLY_ROTARY_POS_EMB_LOOP_6_mux_96_nl
      , APPLY_ROTARY_POS_EMB_LOOP_6_APPLY_ROTARY_POS_EMB_LOOP_6_or_7_nl , APPLY_ROTARY_POS_EMB_LOOP_6_mux_97_nl
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux_98_nl}))) * $signed(({APPLY_ROTARY_POS_EMB_LOOP_6_mux_99_nl
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux_100_nl , APPLY_ROTARY_POS_EMB_LOOP_6_mux_101_nl}));
  assign nl_APPLY_ROTARY_POS_EMB_LOOP_6_mul_sgnd = $signed(({LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48
      , LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_15_8 , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_1 , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_2
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_3 , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_4
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_5 , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_6
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_mux_16_psp_1_ftd_7})) * $signed(({reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd
      , reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1
      , reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2
      , (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3[7:5])
      , 1'b1 , (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3[4:0])}));
  assign nl_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_16_psp_1  = conv_u2u_2_3(TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_15_sdt_1[2:1])
      + conv_u2u_2_3({reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign attention_2_1_16_16_4_4_v_proj_re_mux_nl = MUX_v_24_2_2(output_0_7_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_63_cse);
  assign not_4589_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_44_nl = MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_63_cse);
  assign not_4590_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_36_nl = MUX_v_24_2_2(output_0_8_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_65_cse);
  assign not_4591_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_45_nl = MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_65_cse);
  assign not_4592_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_37_nl = MUX_v_24_2_2(output_0_6_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_67_cse);
  assign not_4593_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_46_nl = MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_67_cse);
  assign not_4594_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_38_nl = MUX_v_24_2_2(output_0_9_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_69_cse);
  assign not_4595_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_47_nl = MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_69_cse);
  assign not_4596_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_39_nl = MUX_v_24_2_2(output_0_5_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_71_cse);
  assign not_4597_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_48_nl = MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_71_cse);
  assign not_4598_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_40_nl = MUX_v_24_2_2(output_0_10_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_73_cse);
  assign not_4599_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_49_nl = MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_73_cse);
  assign not_4600_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_41_nl = MUX_v_24_2_2(output_0_4_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_75_cse);
  assign not_4601_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_50_nl = MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_75_cse);
  assign not_4602_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_42_nl = MUX_v_24_2_2(output_0_11_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_77_cse);
  assign not_4603_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_51_nl = MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_77_cse);
  assign not_4604_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_43_nl = MUX_v_24_2_2(output_0_3_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_79_cse);
  assign not_4605_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_52_nl = MUX_v_16_2_2(apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_79_cse);
  assign not_4606_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_44_nl = MUX_v_24_2_2(output_0_12_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_81_cse);
  assign not_4607_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_53_nl = MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_81_cse);
  assign not_4608_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_45_nl = MUX_v_24_2_2(output_0_2_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_83_cse);
  assign not_4609_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_54_nl = MUX_v_16_2_2(apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_83_cse);
  assign not_4610_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_46_nl = MUX_v_24_2_2(output_0_13_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_85_cse);
  assign not_4611_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_55_nl = MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_85_cse);
  assign not_4612_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_47_nl = MUX_v_24_2_2(output_0_1_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  assign not_4613_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_56_nl = MUX_v_8_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_15_8,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:8]),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  assign not_5055_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_60_nl = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_7,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[7]),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_61_nl = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_6,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[6]),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_62_nl = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_5,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[5]),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_63_nl = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_4,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[4]),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_64_nl = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_3,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[3]),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_65_nl = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_2,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[2]),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_66_nl = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_1,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[1]),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_67_nl = MUX_s_1_2_2(APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_itm_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[0]),
      attention_2_1_16_16_4_4_v_proj_re_and_87_cse);
  assign attention_2_1_16_16_4_4_v_proj_re_mux_48_nl = MUX_v_24_2_2(output_0_14_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_89_cse);
  assign not_4615_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_57_nl = MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_89_cse);
  assign not_4616_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_49_nl = MUX_v_24_2_2(output_0_0_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_91_cse);
  assign not_4617_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_58_nl = MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_91_cse);
  assign not_4618_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_50_nl = MUX_v_24_2_2(output_0_15_sva_1_39_16,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[39:16]),
      attention_2_1_16_16_4_4_v_proj_re_and_93_cse);
  assign not_4619_nl = ~ and_dcpl_1154;
  assign attention_2_1_16_16_4_4_k_proj_re_mux_59_nl = MUX_v_16_2_2(attention_2_1_16_16_4_4_k_proj_2_0_3_lpi_3_15_0,
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_LINEAR_FORWARD_NO_MUL_LOOP_2_2_div_1_cmp_z[15:0]),
      attention_2_1_16_16_4_4_v_proj_re_and_93_cse);
  assign not_4620_nl = ~ and_dcpl_1154;
  assign GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_4_nl = ~(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_5_sva_mx0w0
      & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  assign GEMM_3D_FLOAT_LOOP_3_1_and_32_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_4_nl);
  assign GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_6_nl = ~(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva_mx0w0
      & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  assign GEMM_3D_FLOAT_LOOP_3_1_and_34_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_6_nl);
  assign GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_2_nl = ~(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_6_sva_mx0w0
      & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  assign GEMM_3D_FLOAT_LOOP_3_1_and_30_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_2_nl);
  assign GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_12_nl = ~(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_1_sva_mx0w3
      & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  assign GEMM_3D_FLOAT_LOOP_3_1_and_40_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_12_nl);
  assign GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_10_nl = ~(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva_mx0w3
      & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  assign GEMM_3D_FLOAT_LOOP_3_1_and_38_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_10_nl);
  assign GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_14_nl = ~(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_0_sva_mx0w3
      & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  assign GEMM_3D_FLOAT_LOOP_3_1_and_42_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_14_nl);
  assign mux_789_nl = MUX_s_1_2_2((~ or_tmp_704), and_1651_cse, fsm_output[7]);
  assign and_259_nl = mux_789_nl & and_dcpl_226 & nor_1026_cse & and_dcpl;
  assign and_267_nl = and_dcpl_185 & nor_777_cse & (~ (fsm_output[5])) & and_dcpl_231
      & (fsm_output[7]) & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd) & LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0;
  assign or_1734_nl = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd | (~(LINEAR_FORWARD_NO_MUL_LOOP_4_l_2_0_sva_0
      & (fsm_output[7:6]==2'b11)));
  assign mux_793_nl = MUX_s_1_2_2(mux_792_cse, or_1734_nl, fsm_output[3]);
  assign mux_794_nl = MUX_s_1_2_2(mux_793_nl, or_tmp_708, fsm_output[2]);
  assign nand_307_nl = ~((fsm_output[3]) & (fsm_output[6]) & (fsm_output[7]));
  assign mux_791_nl = MUX_s_1_2_2(or_tmp_708, nand_307_nl, fsm_output[2]);
  assign mux_795_nl = MUX_s_1_2_2(mux_794_nl, mux_791_nl, or_1732_cse);
  assign nand_308_nl = ~(((fsm_output[1]) | (fsm_output[3]) | (fsm_output[6])) &
      (fsm_output[7]));
  assign nand_309_nl = ~(((~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[3])
      | (fsm_output[6])) & (fsm_output[7]));
  assign mux_790_nl = MUX_s_1_2_2(nand_308_nl, nand_309_nl, fsm_output[0]);
  assign mux_796_nl = MUX_s_1_2_2(mux_795_nl, mux_790_nl, fsm_output[4]);
  assign mux_797_nl = MUX_s_1_2_2(mux_796_nl, (~ (fsm_output[7])), fsm_output[5]);
  assign nor_980_nl = ~((fsm_output[1]) | (fsm_output[8]));
  assign nor_981_nl = ~((fsm_output[1]) | (fsm_output[0]) | (fsm_output[8]));
  assign or_1854_nl = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1])
      | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0]);
  assign mux_897_nl = MUX_s_1_2_2(nor_980_nl, nor_981_nl, or_1854_nl);
  assign mux_898_nl = MUX_s_1_2_2(mux_897_nl, (fsm_output[8]), fsm_output[5]);
  assign mux_899_nl = MUX_s_1_2_2(mux_898_nl, nor_tmp_307, fsm_output[3]);
  assign mux_896_nl = MUX_s_1_2_2(nor_tmp_307, (fsm_output[5]), fsm_output[3]);
  assign mux_900_nl = MUX_s_1_2_2(mux_899_nl, mux_896_nl, fsm_output[4]);
  assign or_1857_nl = (fsm_output[6]) | mux_900_nl;
  assign and_380_nl = (fsm_output[5]) & (and_1474_cse | (fsm_output[8]));
  assign mux_894_nl = MUX_s_1_2_2(and_380_nl, or_1851_cse, fsm_output[3]);
  assign mux_895_nl = MUX_s_1_2_2(nor_tmp_307, mux_894_nl, fsm_output[4]);
  assign or_1853_nl = (fsm_output[6]) | mux_895_nl;
  assign mux_901_nl = MUX_s_1_2_2(or_1857_nl, or_1853_nl, fsm_output[2]);
  assign nand_316_nl = ~((fsm_output[3]) & (fsm_output[5]) & (fsm_output[1]) & (~
      (fsm_output[8])));
  assign or_1849_nl = (fsm_output[3]) | (fsm_output[5]) | (~ (fsm_output[1])) | (~
      (fsm_output[0])) | (fsm_output[8]);
  assign mux_891_nl = MUX_s_1_2_2(nand_316_nl, or_1849_nl, fsm_output[4]);
  assign mux_888_nl = MUX_s_1_2_2(or_1848_cse, (fsm_output[8]), fsm_output[5]);
  assign or_1847_nl = nor_305_cse | (fsm_output[8]);
  assign mux_889_nl = MUX_s_1_2_2(mux_888_nl, or_1847_nl, fsm_output[3]);
  assign mux_890_nl = MUX_s_1_2_2(mux_889_nl, (fsm_output[8]), fsm_output[4]);
  assign mux_892_nl = MUX_s_1_2_2(mux_891_nl, mux_890_nl, fsm_output[6]);
  assign or_1846_nl = (~ (fsm_output[4])) | (fsm_output[3]) | (fsm_output[5]) | (fsm_output[1])
      | (fsm_output[0]) | (fsm_output[8]);
  assign or_1845_nl = (~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b00) |
      reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0])
      | (~ (fsm_output[4])) | (fsm_output[3]) | (~ (fsm_output[5])) | (~ (fsm_output[1]))
      | (~ (fsm_output[0])))) | (fsm_output[8]);
  assign mux_887_nl = MUX_s_1_2_2(or_1846_nl, or_1845_nl, fsm_output[6]);
  assign mux_893_nl = MUX_s_1_2_2(mux_892_nl, mux_887_nl, fsm_output[2]);
  assign mux_902_nl = MUX_s_1_2_2(mux_901_nl, mux_893_nl, fsm_output[7]);
  assign GEMM_3D_FLOAT_LOOP_4_1_mux_17_nl = MUX_s_1_16_2((apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2[39]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2[39]), (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2[39]),
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2[39]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2[39]), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2[39]),
      (attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3[39]), (attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3[39]),
      (attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3[39]), (attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3[39]),
      (attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3[39]), (attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3[39]),
      (attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3[39]), (attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3[39]),
      (attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3[39]), {reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign rms_norm_16_variance_mux1h_nl = MUX1HOT_s_1_9_2((acc_3_cse_40_1[39]), (compute_sqrt_for_acc_1_itm_40_1_1[39]),
      attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_39, (APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1[39]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux1h_5_itm[39]), (softmax_1_4_3_sum_sva_2[39]), (SOFTMAX_LOOP_5_mux_12_psp_mx0w0[39]),
      GEMM_3D_FLOAT_LOOP_4_1_mux_17_nl, (compute_sqrt_1_for_acc_1_itm_40_1_1[39]),
      {rms_norm_16_variance_or_1_cse , and_dcpl_290 , and_404_itm , and_dcpl_374
      , and_dcpl_313 , and_dcpl_377 , and_dcpl_294 , and_dcpl_316 , and_dcpl_292});
  assign GEMM_3D_FLOAT_LOOP_4_1_mux_24_nl = MUX_v_39_16_2((apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_2[38:0]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_2[38:0]), (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_2[38:0]),
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_2[38:0]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_2[38:0]), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_2[38:0]),
      (attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3[38:0]), (attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3[38:0]),
      (attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3[38:0]), (attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3[38:0]),
      (attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3[38:0]), (attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3[38:0]),
      (attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3[38:0]), (attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3[38:0]),
      (attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3[38:0]), {reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign rms_norm_16_variance_mux1h_1_nl = MUX1HOT_v_39_10_2((acc_3_cse_40_1[38:0]),
      (compute_sqrt_for_acc_1_itm_40_1_1[38:0]), (attention_abs_1_qr_sva_1[38:0]),
      attention_max_attn_fixed_t_attention_max_attn_fixed_t_and_mut_mx0w3_38_0, (APPLY_ROTARY_POS_EMB_LOOP_3_acc_12_ctmp_sva_1[38:0]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux1h_5_itm[38:0]), (softmax_1_4_3_sum_sva_2[38:0]),
      (SOFTMAX_LOOP_5_mux_12_psp_mx0w0[38:0]), GEMM_3D_FLOAT_LOOP_4_1_mux_24_nl,
      (compute_sqrt_1_for_acc_1_itm_40_1_1[38:0]), {rms_norm_16_variance_or_1_cse
      , and_dcpl_290 , and_dcpl_363 , and_404_itm , and_dcpl_374 , and_dcpl_313 ,
      and_dcpl_377 , and_dcpl_294 , and_dcpl_316 , and_dcpl_292});
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux_nl
      = MUX_s_1_2_2((LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0[3]), (z_out_12[3]),
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_cse);
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_8_nl = MUX1HOT_s_1_5_2((LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0[2]),
      (z_out_12[2]), (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_15_sdt_1[2]), (z_out_3[2]),
      reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1, {and_416_itm , LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_cse
      , LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_7_cse , LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_8_cse
      , LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_9_cse});
  assign and_1238_nl = nor_1314_cse & and_dcpl_200 & and_dcpl_885;
  assign QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux_nl = MUX_v_2_2_2(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2,
      (z_out_3[1:0]), and_1238_nl);
  assign mux_2231_nl = MUX_s_1_2_2((~ nor_tmp_329), or_tmp_1221, fsm_output[3]);
  assign mux_2230_nl = MUX_s_1_2_2(or_tmp_992, or_tmp_861, fsm_output[3]);
  assign mux_2232_nl = MUX_s_1_2_2(mux_2231_nl, mux_2230_nl, fsm_output[6]);
  assign nor_1322_nl = ~(mux_2232_nl | or_1851_cse | (~ (fsm_output[7])));
  assign QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_1_nl
      = MUX_v_2_2_2(2'b00, QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux_nl,
      nor_1322_nl);
  assign nor_996_nl = ~(and_1474_cse | (fsm_output[2]) | (~ (fsm_output[4])));
  assign mux_983_nl = MUX_s_1_2_2(and_1570_cse, nor_996_nl, fsm_output[3]);
  assign mux_982_nl = MUX_s_1_2_2(or_270_cse, or_tmp_861, fsm_output[3]);
  assign mux_984_nl = MUX_s_1_2_2(mux_983_nl, (~ mux_982_nl), fsm_output[6]);
  assign and_426_nl = mux_984_nl & and_dcpl_388;
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_9_nl = MUX1HOT_v_2_6_2((LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0[1:0]),
      (z_out_12[1:0]), QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_1_nl,
      (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_acc_15_sdt_1[1:0]), (z_out_3[1:0]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2,
      {and_416_itm , LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_or_cse , and_426_nl , LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_7_cse
      , LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_8_cse , LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_9_cse});
  assign compute_sqrt_for_i_mux1h_nl = MUX1HOT_s_1_4_2((LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1[3]),
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp[3]), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0[3]),
      (RMS_NORM_LOOP_2_2_i_4_0_sva_1[3]), {and_dcpl_242 , LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c2
      , LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c5 , and_dcpl_410});
  assign compute_sqrt_for_i_mux1h_1_nl = MUX1HOT_v_2_7_2((LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1[2:1]),
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp[2:1]), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0[2:1]),
      (RMS_NORM_LOOP_2_2_i_4_0_sva_1[2:1]), (z_out_5[2:1]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1,
      (z_out_11[2:1]), {and_dcpl_242 , LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c2
      , LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c5 , and_dcpl_410 , compute_sqrt_for_i_and_cse
      , compute_sqrt_for_i_and_4_cse , compute_sqrt_for_i_and_5_cse});
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_not_2_nl = ~ LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c3;
  assign compute_sqrt_for_i_nand_1_nl = ~(MUX_v_2_2_2(2'b00, compute_sqrt_for_i_mux1h_1_nl,
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_not_2_nl));
  assign compute_sqrt_for_i_or_nl = compute_sqrt_for_i_and_4_cse | compute_sqrt_for_i_and_2_cse;
  assign compute_sqrt_for_i_mux1h_2_nl = MUX1HOT_s_1_8_2((LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1[0]),
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp[0]), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0[0]),
      (RMS_NORM_LOOP_2_2_i_4_0_sva_1[0]), (z_out_5[0]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2,
      (z_out_11[0]), (~ QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1),
      {and_dcpl_242 , LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c2 , LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_mx0c5
      , and_dcpl_410 , compute_sqrt_for_i_and_cse , compute_sqrt_for_i_or_nl , compute_sqrt_for_i_and_5_cse
      , and_dcpl_557});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_37_nl = MUX_s_1_16_2(QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39,
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd, (apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_39_16[23]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16[23]), (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3[39]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm[39]), (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_39_16[23]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16[23]), (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3[39]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm[39]), (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_39_16[23]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16[23]), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3[39]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm[39]), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_39_16[23]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16[23]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_69_nl = MUX_v_23_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[38:16]),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1[38:16]), (apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_39_16[22:0]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16[22:0]), (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3[38:16]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm[38:16]), (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_39_16[22:0]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16[22:0]), (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3[38:16]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm[38:16]), (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_39_16[22:0]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_39_16[22:0]), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3[38:16]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm[38:16]), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_39_16[22:0]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_39_16[22:0]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign nand_373_nl = ~((reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0 | (~ reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1)
      | reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 | reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd)
      & (fsm_output[2]) & (fsm_output[3]) & (fsm_output[1]) & (fsm_output[0]) & (~
      (fsm_output[6])) & (fsm_output[7]));
  assign nor_576_nl = ~((~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      | (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1))) | (fsm_output[3:0]!=4'b0001));
  assign mux_2079_nl = MUX_s_1_2_2(or_1983_cse, mux_806_cse, nor_576_nl);
  assign mux_2080_nl = MUX_s_1_2_2(nand_373_nl, mux_2079_nl, fsm_output[4]);
  assign or_2775_nl = (fsm_output[1]) | (fsm_output[0]) | (~ (fsm_output[6])) | (fsm_output[7]);
  assign mux_2077_nl = MUX_s_1_2_2(or_1983_cse, or_2775_nl, and_1773_cse);
  assign or_2777_nl = (fsm_output[4]) | mux_2077_nl;
  assign mux_2081_nl = MUX_s_1_2_2(mux_2080_nl, or_2777_nl, fsm_output[5]);
  assign nor_1225_nl = ~(mux_2081_nl | (fsm_output[8]));
  assign and_1110_nl = and_dcpl_1061 & and_dcpl_45 & (~ reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd)
      & (~(reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1 | reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0))
      & reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1;
  assign and_1115_nl = and_dcpl_205 & and_dcpl_421 & and_dcpl_319 & (~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd)) & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign INIT_2D_MEM_LOOP_2_1_mux1h_nl = MUX1HOT_v_24_9_2(attention_2_1_16_16_4_4_v_proj_re_0_10_sva_1_39_16,
      LINEAR_FORWARD_NO_MUL_LOOP_2_2_conc_1_mut_71_48_mx0w0, for_for_strm_in_tmp_sva_25_2,
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_39_16,
      RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_39_16, APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1,
      ({APPLY_ROTARY_POS_EMB_LOOP_6_mux_37_nl , APPLY_ROTARY_POS_EMB_LOOP_6_mux_69_nl}),
      {and_dcpl_726 , and_dcpl_257 , nor_1225_nl , and_dcpl_1011 , and_dcpl_983 ,
      and_1110_nl , and_dcpl_847 , and_1115_nl , and_dcpl_583});
  assign mux_2074_nl = MUX_s_1_2_2((~ or_tmp_728), or_tmp_767, fsm_output[5]);
  assign mux_2075_nl = MUX_s_1_2_2(mux_tmp_91, mux_2074_nl, fsm_output[3]);
  assign nand_96_nl = ~((fsm_output[6]) & (~ mux_2075_nl));
  assign mux_2076_nl = MUX_s_1_2_2(nand_96_nl, or_tmp_913, fsm_output[7]);
  assign nor_1323_nl = ~(mux_2076_nl | (fsm_output[8]));
  assign INIT_2D_MEM_LOOP_2_1_and_nl = MUX_v_24_2_2(24'b000000000000000000000000,
      INIT_2D_MEM_LOOP_2_1_mux1h_nl, nor_1323_nl);
  assign GEMM_3D_FLOAT_LOOP_4_mux_17_nl = MUX_v_40_16_2(attention_2_1_16_16_4_4_q_embed_0_0_0_sva_1,
      attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1, attention_2_1_16_16_4_4_q_embed_0_0_2_sva_1,
      attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1, attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1,
      attention_2_1_16_16_4_4_q_embed_1_0_1_sva_1, attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1,
      attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1, attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1,
      attention_2_1_16_16_4_4_q_embed_2_0_1_sva_1, attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1,
      attention_2_1_16_16_4_4_q_embed_2_0_3_sva_1, attention_2_1_16_16_4_4_q_embed_3_0_0_sva_1,
      attention_2_1_16_16_4_4_q_embed_3_0_1_sva_1, attention_2_1_16_16_4_4_q_embed_3_0_2_sva_1,
      attention_2_1_16_16_4_4_q_embed_3_0_3_sva_1, {reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1});
  assign SOFTMAX_LOOP_4_x_mux_nl = MUX_v_40_12_2(attention_2_1_16_16_4_4_attn_weights_0_0_0_lpi_9,
      attention_2_1_16_16_4_4_attn_weights_1_0_0_lpi_9, attention_2_1_16_16_4_4_attn_weights_2_0_0_lpi_9,
      attention_2_1_16_16_4_4_attn_weights_3_0_0_lpi_9, attention_2_1_16_16_4_4_attn_weights_0_0_1_lpi_8,
      attention_2_1_16_16_4_4_attn_weights_1_0_1_lpi_8, attention_2_1_16_16_4_4_attn_weights_2_0_1_lpi_8,
      attention_2_1_16_16_4_4_attn_weights_3_0_1_lpi_8, attention_2_1_16_16_4_4_attn_weights_0_0_2_lpi_8,
      attention_2_1_16_16_4_4_attn_weights_1_0_2_lpi_8, attention_2_1_16_16_4_4_attn_weights_2_0_2_lpi_8,
      attention_2_1_16_16_4_4_attn_weights_3_0_2_lpi_8, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign nl_SOFTMAX_LOOP_4_x_acc_2_nl = SOFTMAX_LOOP_4_x_mux_nl + ({(~ QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39)
      , (~ QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0)}) + 40'b0000000000000000000000000000000000000001;
  assign SOFTMAX_LOOP_4_x_acc_2_nl = nl_SOFTMAX_LOOP_4_x_acc_2_nl[39:0];
  assign GEMM_3D_FLOAT_LOOP_4_1_mux_18_nl = MUX_v_40_12_2(attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1, {reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2
      , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd , reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign mux_1059_nl = MUX_s_1_2_2(or_tmp_930, mux_tmp_1044, fsm_output[1]);
  assign mux_1058_nl = MUX_s_1_2_2(or_tmp_930, or_tmp_931, fsm_output[1]);
  assign mux_1060_nl = MUX_s_1_2_2(mux_1059_nl, mux_1058_nl, fsm_output[0]);
  assign mux_1057_nl = MUX_s_1_2_2(mux_tmp_1051, or_tmp_930, fsm_output[1]);
  assign mux_1061_nl = MUX_s_1_2_2(mux_1060_nl, mux_1057_nl, fsm_output[3]);
  assign mux_1054_nl = MUX_s_1_2_2(or_tmp_931, mux_tmp_1052, fsm_output[1]);
  assign mux_1053_nl = MUX_s_1_2_2(mux_tmp_1052, mux_tmp_1051, fsm_output[1]);
  assign mux_1055_nl = MUX_s_1_2_2(mux_1054_nl, mux_1053_nl, fsm_output[0]);
  assign or_1996_nl = (fsm_output[1]) | (fsm_output[4]) | (~ (fsm_output[7]));
  assign mux_1050_nl = MUX_s_1_2_2(or_tmp_930, or_1996_nl, fsm_output[0]);
  assign mux_1056_nl = MUX_s_1_2_2(mux_1055_nl, mux_1050_nl, fsm_output[3]);
  assign mux_1062_nl = MUX_s_1_2_2(mux_1061_nl, mux_1056_nl, fsm_output[2]);
  assign or_1994_nl = nor_646_cse | (fsm_output[7]);
  assign mux_1047_nl = MUX_s_1_2_2((~ mux_tmp_1044), (fsm_output[7]), or_1732_cse);
  assign mux_1048_nl = MUX_s_1_2_2(or_1994_nl, mux_1047_nl, fsm_output[3]);
  assign mux_1042_nl = MUX_s_1_2_2((fsm_output[7]), (~ (fsm_output[7])), fsm_output[4]);
  assign mux_1043_nl = MUX_s_1_2_2(mux_1042_nl, or_tmp_922, fsm_output[5]);
  assign mux_1045_nl = MUX_s_1_2_2(mux_tmp_1044, mux_1043_nl, nor_366_cse);
  assign mux_1046_nl = MUX_s_1_2_2((~ mux_1045_nl), (fsm_output[7]), fsm_output[3]);
  assign mux_1049_nl = MUX_s_1_2_2(mux_1048_nl, mux_1046_nl, fsm_output[2]);
  assign mux_1063_nl = MUX_s_1_2_2(mux_1062_nl, mux_1049_nl, fsm_output[6]);
  assign RMS_NORM_LOOP_2_mux_22_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1[39]),
      (input_0_1_sva_1[39]), input_0_2_sva_1_39, (input_0_3_sva_1[39]), (input_0_4_sva_1[39]),
      (input_0_5_sva_1[39]), (input_0_6_sva_1[39]), (input_0_7_sva_1[39]), (input_0_8_sva_1[39]),
      (input_0_9_sva_1[39]), (input_0_10_sva_1[39]), (input_0_11_sva_1[39]), (input_0_12_sva_1[39]),
      input_0_13_sva_1_39, (input_0_14_sva_1[39]), (attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3[39]),
      {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
  assign QUANTIZE_ACTIVATION_LOOP_3_quantized_value_mux_nl = MUX_s_1_16_2((input_0_0_sva_2[39]),
      (input_0_1_sva_2[39]), input_0_2_sva_2_39, (input_0_3_sva_2[39]), (input_0_4_sva_2[39]),
      (input_0_5_sva_2[39]), (input_0_6_sva_2[39]), (input_0_7_sva_2[39]), (input_0_8_sva_2[39]),
      (input_0_9_sva_2[39]), (input_0_10_sva_2[39]), (input_0_11_sva_2[39]), (input_0_12_sva_2[39]),
      input_0_13_sva_2_39, (input_0_14_sva_2[39]), (input_0_15_sva_1[39]), {reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2});
  assign RMS_NORM_LOOP_2_mux_24_nl = MUX_v_39_16_2((attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1[38:0]),
      (input_0_1_sva_1[38:0]), input_0_2_sva_1_38_0, (input_0_3_sva_1[38:0]), (input_0_4_sva_1[38:0]),
      (input_0_5_sva_1[38:0]), (input_0_6_sva_1[38:0]), (input_0_7_sva_1[38:0]),
      (input_0_8_sva_1[38:0]), (input_0_9_sva_1[38:0]), (input_0_10_sva_1[38:0]),
      (input_0_11_sva_1[38:0]), (input_0_12_sva_1[38:0]), input_0_13_sva_1_38_0,
      (input_0_14_sva_1[38:0]), (attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3[38:0]),
      {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
  assign QUANTIZE_ACTIVATION_LOOP_3_quantized_value_mux_1_nl = MUX_v_39_16_2((input_0_0_sva_2[38:0]),
      (input_0_1_sva_2[38:0]), input_0_2_sva_2_38_0, (input_0_3_sva_2[38:0]), (input_0_4_sva_2[38:0]),
      (input_0_5_sva_2[38:0]), (input_0_6_sva_2[38:0]), (input_0_7_sva_2[38:0]),
      (input_0_8_sva_2[38:0]), (input_0_9_sva_2[38:0]), (input_0_10_sva_2[38:0]),
      (input_0_11_sva_2[38:0]), (input_0_12_sva_2[38:0]), input_0_13_sva_2_38_0,
      (input_0_14_sva_2[38:0]), (input_0_15_sva_1[38:0]), {reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1 , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2});
  assign for_for_for_for_nand_nl = ~(mux_1079_itm & (~(or_dcpl_1025 & and_dcpl_204)));
  assign for_for_and_24_nl = (~ or_dcpl_1025) & and_dcpl_204;
  assign for_for_mux1h_5_nl = MUX1HOT_v_40_9_2(({{10{strm_in_rsci_idat_mxwt[29]}},
      strm_in_rsci_idat_mxwt}), input_0_12_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1, attention_2_1_16_16_4_4_q_embed_0_0_0_sva_1,
      attention_2_1_16_16_4_4_attn_weights_1_0_0_sva_2, attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx2,
      ({ATTN_2D_LOOP_3_mux_16_itm , ATTN_2D_LOOP_3_mux_17_itm}), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      {attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c0 , attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c1
      , for_for_for_for_nand_nl , for_for_and_24_nl , and_dcpl_216 , and_dcpl_348
      , and_dcpl_351 , and_dcpl_352 , attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c9});
  assign attention_2_1_16_16_4_4_attn_output_2D_not_nl = ~ attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1_mx0c7;
  assign for_for_mux1h_6_nl = MUX1HOT_v_40_8_2(({{10{strm_in_rsci_idat_mxwt[29]}},
      strm_in_rsci_idat_mxwt}), input_0_7_sva_1, attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1,
      attention_2_1_16_16_4_4_q_embed_0_0_1_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_weights_2_0_2_sva_2,
      attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx1, ({ATTN_2D_LOOP_3_mux_16_itm
      , ATTN_2D_LOOP_3_mux_17_itm}), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      {attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c0 , attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c1
      , and_dcpl_346 , and_dcpl_204 , and_dcpl_348 , and_dcpl_351 , and_dcpl_352
      , attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c9});
  assign attention_2_1_16_16_4_4_attn_output_2D_not_3_nl = ~ attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1_mx0c7;
  assign or_2048_nl = (~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b10) |
      reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 | (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]))
      | (fsm_output[4:0]!=5'b10111))) | (fsm_output[8]);
  assign mux_1095_nl = MUX_s_1_2_2(mux_1074_cse, or_2048_nl, fsm_output[5]);
  assign mux_1097_nl = MUX_s_1_2_2(nand_50_cse, mux_1095_nl, fsm_output[6]);
  assign mux_1099_nl = MUX_s_1_2_2(or_2029_cse, mux_1097_nl, fsm_output[7]);
  assign GEMM_3D_FLOAT_LOOP_3_1_and_36_nl = reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd
      & GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_8_seb;
  assign GEMM_3D_FLOAT_LOOP_3_1_and_52_nl = MUX_v_39_2_2(39'b000000000000000000000000000000000000000,
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_8_seb);
  assign for_for_and_22_nl = (~ and_dcpl_548) & and_dcpl_477;
  assign GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_nl = ~(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_7_sva_mx0w0
      & (~ reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd));
  assign GEMM_3D_FLOAT_LOOP_3_1_and_28_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_1_0_3_lpi_3, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_nl);
  assign and_521_nl = and_dcpl_342 & and_dcpl_336 & and_dcpl_480;
  assign and_523_nl = or_dcpl_1084 & and_dcpl_185 & and_dcpl_422;
  assign GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_1_nl = ~(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_0_sva_mx0w3
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd);
  assign GEMM_3D_FLOAT_LOOP_3_1_and_29_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2_0_0_lpi_3, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_1_nl);
  assign and_527_nl = and_dcpl_342 & and_dcpl_417 & and_dcpl_486;
  assign and_529_nl = or_dcpl_1085 & and_dcpl_185 & and_dcpl_422;
  assign GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_3_nl = ~(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_1_sva_mx0w3
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd);
  assign GEMM_3D_FLOAT_LOOP_3_1_and_31_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2_0_1_lpi_3, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_3_nl);
  assign and_531_nl = and_dcpl_342 & and_dcpl_336 & and_dcpl_486;
  assign and_533_nl = or_dcpl_1086 & and_dcpl_185 & and_dcpl_422;
  assign GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_5_nl = ~(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_2_sva_mx0w3
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd);
  assign GEMM_3D_FLOAT_LOOP_3_1_and_33_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2_0_2_lpi_3, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_5_nl);
  assign and_535_nl = and_dcpl_342 & and_dcpl_417 & and_dcpl_480;
  assign and_537_nl = or_dcpl_1087 & and_dcpl_185 & and_dcpl_422;
  assign GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_7_nl = ~(GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_3_sva_mx0w3
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd);
  assign GEMM_3D_FLOAT_LOOP_3_1_and_35_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2_0_3_lpi_3, GEMM_3D_FLOAT_LOOP_3_1_GEMM_3D_FLOAT_LOOP_3_1_nand_7_nl);
  assign and_539_nl = and_dcpl_342 & and_dcpl_336 & and_dcpl_471;
  assign and_541_nl = or_dcpl_1088 & and_dcpl_185 & and_dcpl_422;
  assign for_for_or_4_nl = attention_2_1_16_16_4_4_q_embed_and_24_cse | and_dcpl_222
      | (nand_302_cse & and_dcpl_187);
  assign for_for_and_28_nl = (~ nand_302_cse) & and_dcpl_187;
  assign for_for_mux1h_13_nl = MUX1HOT_v_40_8_2(({{10{strm_in_rsci_idat_mxwt[29]}},
      strm_in_rsci_idat_mxwt}), input_0_10_sva_1, attention_2_1_16_16_4_4_k_embed_2_0_3_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1, attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3,
      acc_3_cse_40_1, ({ATTN_2D_LOOP_3_mux_16_itm , ATTN_2D_LOOP_3_mux_17_itm}),
      RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva, {attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c0
      , attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c1 , and_dcpl_346 , attention_2_1_16_16_4_4_q_embed_and_23_cse
      , for_for_or_4_nl , for_for_and_28_nl , and_dcpl_352 , attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c10});
  assign for_for_or_3_nl = MUX_v_40_2_2(for_for_mux1h_13_nl, 40'b1111111111111111111111111111111111111111,
      attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c8);
  assign or_nl = ((~ (z_out_5[2])) & attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c8)
      | attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c5;
  assign mux_nl = MUX_v_40_2_2(for_for_or_3_nl, attention_2_1_16_16_4_4_attn_output_3_0_0_sva_2,
      or_nl);
  assign nor_nl = ~((GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_4_sva_mx0w0 & and_dcpl_222
      & reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd) | ((z_out_5[2]) & attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3_mx0c8));
  assign or_2087_nl = (~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b11) |
      reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0])
      | (fsm_output[4:0]!=5'b10111))) | (fsm_output[8:6]!=3'b011);
  assign mux_1133_nl = MUX_s_1_2_2(mux_1132_cse, or_2087_nl, fsm_output[5]);
  assign or_3215_nl = (~ mux_1147_itm) | (and_dcpl_222 & (~ or_3212_tmp)) | attention_2_1_16_16_4_4_attn_output_and_14_cse
      | attention_2_1_16_16_4_4_q_embed_and_26_cse;
  assign mux1h_nl = MUX1HOT_v_40_9_2(({{10{strm_in_rsci_idat_mxwt[29]}}, strm_in_rsci_idat_mxwt}),
      input_0_4_sva_1, attention_2_1_16_16_4_4_k_embed_3_0_0_sva_1, attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1, attention_2_1_16_16_4_4_attn_output_3_0_1_sva_2,
      acc_3_cse_40_1, ({ATTN_2D_LOOP_3_mux_16_itm , ATTN_2D_LOOP_3_mux_17_itm}),
      RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva, {attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c0
      , attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c1 , and_dcpl_346 , or_3215_nl
      , attention_2_1_16_16_4_4_q_embed_and_25_cse , and_dcpl_524 , attention_2_1_16_16_4_4_attn_output_and_13_cse
      , and_dcpl_352 , attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3_mx0c10});
  assign not_4622_nl = ~ or_3212_tmp;
  assign or_3216_nl = (~ mux_1177_itm) | (and_dcpl_222 & (~ or_3213_tmp)) | attention_2_1_16_16_4_4_attn_output_and_16_cse
      | attention_2_1_16_16_4_4_q_embed_and_28_cse;
  assign mux1h_1_nl = MUX1HOT_v_40_9_2(({{10{strm_in_rsci_idat_mxwt[29]}}, strm_in_rsci_idat_mxwt}),
      input_0_11_sva_1, attention_2_1_16_16_4_4_k_embed_3_0_1_sva_1, attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1, attention_2_1_16_16_4_4_attn_output_3_0_2_sva_2,
      acc_3_cse_40_1, ({ATTN_2D_LOOP_3_mux_16_itm , ATTN_2D_LOOP_3_mux_17_itm}),
      RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva, {attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c0
      , attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c1 , and_dcpl_346 , or_3216_nl
      , attention_2_1_16_16_4_4_q_embed_and_27_cse , and_dcpl_524 , attention_2_1_16_16_4_4_attn_output_and_15_cse
      , and_dcpl_352 , attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3_mx0c10});
  assign not_4624_nl = ~ or_3213_tmp;
  assign or_3217_nl = (~ mux_1197_itm) | (and_dcpl_222 & (~ or_3214_tmp)) | attention_2_1_16_16_4_4_attn_output_and_18_cse
      | attention_2_1_16_16_4_4_q_embed_and_30_cse;
  assign mux1h_2_nl = MUX1HOT_v_40_11_2(({{10{strm_in_rsci_idat_mxwt[29]}}, strm_in_rsci_idat_mxwt}),
      input_0_3_sva_1, (signext_40_30({for_for_strm_in_tmp_sva_31_26 , for_for_strm_in_tmp_sva_25_2})),
      attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3, input_0_15_sva_1, attention_2_1_16_16_4_4_k_embed_3_0_2_sva_1,
      APPLY_ROTARY_POS_EMB_LOOP_6_acc_14_itm_55_16_1, attention_2_1_16_16_4_4_attn_output_3_0_3_sva_2,
      acc_3_cse_40_1, ({ATTN_2D_LOOP_3_mux_16_itm , ATTN_2D_LOOP_3_mux_17_itm}),
      RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva, {attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c0
      , attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c1 , and_dcpl_242 , or_3217_nl
      , and_dcpl_344 , and_dcpl_346 , attention_2_1_16_16_4_4_q_embed_and_29_cse
      , and_dcpl_524 , attention_2_1_16_16_4_4_attn_output_and_17_cse , and_dcpl_352
      , attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3_mx0c12});
  assign not_4626_nl = ~ or_3214_tmp;
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_7_nl = MUX1HOT_s_1_5_2((z_out_12[4]),
      (compute_sqrt_for_acc_1_itm_40_1_1[39]), (LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp[4]),
      (compute_sqrt_1_for_acc_1_itm_40_1_1[39]), (RMS_NORM_LOOP_2_2_acc_1_tmp[4]),
      {and_581_ssc , and_dcpl_290 , and_dcpl_439 , and_dcpl_292 , and_dcpl_306});
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_10_nl = MUX1HOT_v_4_6_2((z_out_12[3:0]),
      (compute_sqrt_for_acc_1_itm_40_1_1[38:35]), ({reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2}),
      (LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp[3:0]), (compute_sqrt_1_for_acc_1_itm_40_1_1[38:35]),
      (RMS_NORM_LOOP_2_2_acc_1_tmp[3:0]), {and_581_ssc , and_dcpl_290 , and_dcpl_477
      , and_dcpl_439 , and_dcpl_292 , and_dcpl_306});
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_and_4_nl = MUX_v_4_2_2(4'b0000, LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_mux1h_10_nl,
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_nand_seb);
  assign attention_2_1_16_16_4_4_q_proj_attention_2_1_16_16_4_4_q_proj_mux_12_nl
      = MUX_s_1_2_2(attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_15, (z_out[15]), and_1191_rgt);
  assign operator_40_24_true_AC_TRN_AC_WRAP_1_and_2_nl = (~ and_dcpl_739) & (~ mux_1309_cse)
      & (fsm_output[2]) & and_dcpl_577 & and_dcpl_576;
  assign RMS_NORM_LOOP_2_2_i_mux1h_3_nl = MUX1HOT_v_3_3_2((RMS_NORM_LOOP_2_2_i_4_0_sva_1[3:1]),
      (LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1[3:1]), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0[3:1]),
      {and_dcpl_477 , and_dcpl_410 , and_dcpl_255});
  assign RMS_NORM_LOOP_2_2_i_not_2_nl = ~ RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_mx0c1;
  assign APPLY_ROTARY_POS_EMB_LOOP_3_and_10_nl = reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      & (~ reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1);
  assign RMS_NORM_LOOP_2_2_i_mux1h_6_nl = MUX1HOT_s_1_7_2((RMS_NORM_LOOP_2_2_i_4_0_sva_1[0]),
      (LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1[0]), APPLY_ROTARY_POS_EMB_LOOP_3_and_10_nl,
      GEMM_3D_FLOAT_LOOP_3_and_tmp_5_sva_mx0w2, GEMM_3D_FLOAT_LOOP_3_1_and_stg_2_1_sva_mx0w3,
      (~ QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1), (LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0[0]),
      {and_dcpl_477 , and_dcpl_410 , RMS_NORM_LOOP_2_2_i_and_9_cse , and_dcpl_1152
      , and_dcpl_222 , and_dcpl_557 , and_dcpl_255});
  assign or_2335_nl = and_1638_cse | (fsm_output[7:6]!=2'b10);
  assign mux_1433_nl = MUX_s_1_2_2(or_2335_nl, or_1983_cse, fsm_output[5]);
  assign mux_1428_nl = MUX_s_1_2_2(or_1983_cse, (~ (fsm_output[6])), fsm_output[0]);
  assign nor_1105_nl = ~((fsm_output[7:6]!=2'b10));
  assign mux_1429_nl = MUX_s_1_2_2(mux_1428_nl, nor_1105_nl, fsm_output[1]);
  assign mux_1430_nl = MUX_s_1_2_2(or_1983_cse, mux_1429_nl, fsm_output[2]);
  assign or_2331_nl = (~(nor_1106_cse | (fsm_output[6]))) | (fsm_output[7]);
  assign mux_1431_nl = MUX_s_1_2_2(mux_1430_nl, or_2331_nl, fsm_output[3]);
  assign mux_1432_nl = MUX_s_1_2_2(or_1983_cse, mux_1431_nl, fsm_output[5]);
  assign mux_1434_nl = MUX_s_1_2_2(mux_1433_nl, mux_1432_nl, fsm_output[4]);
  assign QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_nl = MUX1HOT_s_1_3_2(reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0,
      (z_out_3[1]), (z_out_3[1]), {QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_or_cse
      , and_dcpl_726 , and_937_ssc});
  assign QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_3_nl = QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_nl
      & nor_1324_seb;
  assign RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_and_nl = (LINEAR_FORWARD_NO_MUL_LOOP_2_2_acc_2_tmp[4])
      & RMS_NORM_LOOP_2_2_unequal_tmp_mx0w0;
  assign QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_3_nl = MUX1HOT_s_1_3_2(reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1,
      (z_out_3[0]), (z_out_3[0]), {QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_or_cse
      , and_dcpl_726 , and_937_ssc});
  assign QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_and_4_nl = QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_qif_mux1h_3_nl
      & nor_1324_seb;
  assign nor_1109_nl = ~((fsm_output[6]) | mux_tmp_1440);
  assign nor_1110_nl = ~((~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2])));
  assign mux_1441_nl = MUX_s_1_2_2(nor_1109_nl, nor_1110_nl, fsm_output[7]);
  assign CACHE_UPDATE_LOOP_3_k_and_1_nl = (~ and_dcpl_629) & mux_1441_nl & and_dcpl_628;
  assign or_594_nl = reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 | reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1;
  assign RMS_NORM_LOOP_2_2_mux1h_nl = MUX1HOT_s_1_3_2(RMS_NORM_LOOP_2_2_unequal_tmp_mx0w0,
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1, or_594_nl, {and_dcpl_386 , and_dcpl_629
      , and_dcpl_207});
  assign nand_348_nl = ~((fsm_output[5]) & and_1637_cse);
  assign or_2341_nl = (~ (fsm_output[5])) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[2]);
  assign mux_1438_nl = MUX_s_1_2_2(nand_348_nl, or_2341_nl, fsm_output[3]);
  assign or_2342_nl = (fsm_output[6]) | mux_1438_nl;
  assign or_2340_nl = (fsm_output[3]) | (fsm_output[5]) | (~ (fsm_output[0])) | (fsm_output[1])
      | (fsm_output[2]);
  assign or_2339_nl = (fsm_output[3]) | (~((fsm_output[5]) & (fsm_output[2])));
  assign mux_1437_nl = MUX_s_1_2_2(or_2340_nl, or_2339_nl, fsm_output[6]);
  assign mux_1439_nl = MUX_s_1_2_2(or_2342_nl, mux_1437_nl, fsm_output[7]);
  assign RMS_NORM_LOOP_2_2_and_36_nl = RMS_NORM_LOOP_2_2_mux1h_nl & (~(mux_1439_nl
      | or_tmp_48));
  assign GEMM_3D_FLOAT_LOOP_1_i_mux_1_nl = MUX_s_1_2_2(RMS_NORM_LOOP_2_2_and_36_nl,
      (z_out_5[0]), GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_mx0c1);
  assign and_688_nl = or_dcpl_1108 & and_dcpl_202 & and_dcpl_642;
  assign and_693_nl = or_dcpl_1114 & and_dcpl_202 & and_dcpl_642;
  assign and_704_nl = or_dcpl_1118 & and_dcpl_202 & and_dcpl_642;
  assign and_709_nl = or_dcpl_1120 & and_dcpl_202 & and_dcpl_642;
  assign and_713_nl = or_dcpl_1121 & and_dcpl_202 & and_dcpl_642;
  assign and_717_nl = or_dcpl_1122 & and_dcpl_202 & and_dcpl_642;
  assign and_721_nl = or_dcpl_1123 & and_dcpl_202 & and_dcpl_642;
  assign and_725_nl = or_dcpl_1125 & and_dcpl_202 & and_dcpl_642;
  assign and_729_nl = or_dcpl_1126 & and_dcpl_202 & and_dcpl_642;
  assign and_733_nl = or_dcpl_1127 & and_dcpl_202 & and_dcpl_642;
  assign and_737_nl = or_dcpl_1128 & and_dcpl_202 & and_dcpl_642;
  assign and_741_nl = or_dcpl_1130 & and_dcpl_202 & and_dcpl_642;
  assign and_749_nl = or_dcpl_1132 & and_dcpl_202 & and_dcpl_642;
  assign and_753_nl = or_dcpl_1133 & and_dcpl_202 & and_dcpl_642;
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_and_1_nl = (LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1[4])
      & LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_4 & (RMS_NORM_LOOP_2_2_i_4_0_sva_1[4]);
  assign and_755_nl = and_dcpl_215 & nor_1138_m1c;
  assign nand_353_nl = ~((fsm_output[6:0]==7'b1111111));
  assign mux_1491_nl = MUX_s_1_2_2(nand_353_nl, or_tmp_1218, fsm_output[7]);
  assign nor_1136_nl = ~(mux_1491_nl | (fsm_output[8]));
  assign and_757_nl = and_dcpl_291 & nor_1138_m1c;
  assign nand_356_nl = ~((fsm_output[5]) & (fsm_output[0]) & (fsm_output[2]) & (~
      (fsm_output[4])));
  assign mux_1514_nl = MUX_s_1_2_2((~ and_1570_cse), or_tmp_1221, fsm_output[0]);
  assign mux_1515_nl = MUX_s_1_2_2(mux_1514_nl, mux_1513_cse, fsm_output[5]);
  assign mux_1516_nl = MUX_s_1_2_2(nand_356_nl, mux_1515_nl, fsm_output[3]);
  assign nor_1141_nl = ~(RESHAPE_2D_TO_3D_LOOP_2_2_and_cse | (fsm_output[3]) | (~
      (fsm_output[4])) | (fsm_output[6]));
  assign nor_1142_nl = ~((fsm_output[1]) | (~ (fsm_output[3])) | (fsm_output[4])
      | (~ (fsm_output[6])));
  assign mux_1536_nl = MUX_s_1_2_2(nor_1141_nl, nor_1142_nl, fsm_output[0]);
  assign or_2463_nl = (~ (fsm_output[3])) | (fsm_output[4]) | (~ (fsm_output[6]));
  assign or_2461_nl = (z_out_4[2]) | (fsm_output[3]) | (~ (fsm_output[4])) | (fsm_output[6]);
  assign mux_1534_nl = MUX_s_1_2_2(or_2463_nl, or_2461_nl, fsm_output[1]);
  assign nor_1143_nl = ~((fsm_output[0]) | mux_1534_nl);
  assign mux_1537_nl = MUX_s_1_2_2(mux_1536_nl, nor_1143_nl, fsm_output[2]);
  assign APPLY_ROTARY_POS_EMB_LOOP_1_i_or_nl = ((~ mux_1309_cse) & and_1559_cse &
      nor_1026_cse & and_dcpl_576) | ((~ mux_1516_nl) & and_dcpl_718) | (mux_1537_nl
      & and_dcpl_388);
  assign APPLY_ROTARY_POS_EMB_LOOP_1_i_mux1h_5_nl = MUX1HOT_s_1_5_2(and_28_cse, LINEAR_FORWARD_NO_MUL_LOOP_2_and_1_nl,
      reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1, RMS_NORM_LOOP_2_2_and_32_ssc_mx0w3,
      (z_out_4[0]), {and_dcpl_363 , and_755_nl , nor_1136_nl , and_757_nl , APPLY_ROTARY_POS_EMB_LOOP_1_i_or_nl});
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_4_nl = MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_v_proj_re_0_15_lpi_4_39_16_mx1,
      attention_2_1_16_16_4_4_v_proj_re_0_15_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_39_16,
      {and_dcpl_725 , and_dcpl_726 , and_dcpl_410});
  assign not_4557_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_8_nl = MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_v_proj_re_0_0_lpi_4_39_16_mx1,
      attention_2_1_16_16_4_4_v_proj_re_0_0_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_39_16,
      {and_dcpl_725 , and_dcpl_726 , and_dcpl_410});
  assign not_4558_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_12_nl = MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_v_proj_re_0_1_lpi_4_39_16_mx1,
      attention_2_1_16_16_4_4_v_proj_re_0_1_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_39_16,
      {and_dcpl_725 , and_dcpl_726 , and_dcpl_410});
  assign not_4559_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_16_nl = MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_v_proj_re_0_3_lpi_4_39_16_mx1,
      attention_2_1_16_16_4_4_v_proj_re_0_3_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_39_16,
      {and_dcpl_725 , and_dcpl_726 , and_dcpl_410});
  assign not_4560_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_20_nl = MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_v_proj_re_0_7_lpi_4_39_16_mx1,
      attention_2_1_16_16_4_4_v_proj_re_0_7_sva_1_39_16, attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_39_16,
      {and_dcpl_725 , and_dcpl_726 , and_dcpl_410});
  assign not_4561_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_21_nl = MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_39_16_mx1,
      attention_2_1_16_16_4_4_k_proj_re_0_7_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_re_0_7_sva_2_39_16,
      {and_dcpl_725 , and_dcpl_726 , and_dcpl_410});
  assign not_4562_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_35_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_7_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_754);
  assign not_4441_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_34_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_8_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_760);
  assign not_4440_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_33_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_6_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_764);
  assign not_4439_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_32_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_9_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_768);
  assign not_4438_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_31_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_5_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_772);
  assign not_4437_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_30_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_10_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_776);
  assign not_4436_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_29_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_4_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_780);
  assign not_4435_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_28_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_11_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_784);
  assign not_4434_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_27_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_12_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_788);
  assign not_4433_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_26_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_13_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_792);
  assign not_4432_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_25_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_1_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_796);
  assign not_4431_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_24_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_14_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_800);
  assign not_4430_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_23_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_0_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_804);
  assign not_4429_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_22_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_q_proj_re_0_15_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_812);
  assign not_4428_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_21_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_8_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_821);
  assign not_4427_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_20_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_6_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_827);
  assign not_4426_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_19_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_9_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_832);
  assign not_4425_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_18_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_5_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_837);
  assign not_4424_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_17_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_4_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_851);
  assign not_4422_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux_16_nl = MUX_v_24_2_2(attention_2_1_16_16_4_4_k_proj_re_0_15_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), and_dcpl_880);
  assign not_4415_nl = ~ and_dcpl_619;
  assign and_1184_nl = or_dcpl_1141 & and_dcpl_191 & and_dcpl_641 & and_dcpl_813;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_40_nl = MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_re_0_10_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_2_0_3_sva_1_39_16, {attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_3_39_16_mx0c1
      , and_dcpl_843 , and_dcpl_207 , and_dcpl_847});
  assign not_4423_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_42_nl = MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_re_0_11_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_3_0_0_sva_1_39_16, {attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_3_39_16_mx0c1
      , and_dcpl_856 , and_dcpl_207 , and_dcpl_847});
  assign not_4421_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_43_nl = MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_re_0_12_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_3_0_1_sva_1_39_16, {attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_3_39_16_mx0c1
      , and_dcpl_860 , and_dcpl_207 , and_dcpl_847});
  assign not_4420_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_44_nl = MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_re_0_13_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_3_0_2_sva_1_39_16, {attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_3_39_16_mx0c1
      , and_dcpl_864 , and_dcpl_207 , and_dcpl_847});
  assign not_4419_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_45_nl = MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_re_0_1_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_2_0_2_sva_1_39_16, {attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_3_39_16_mx0c1
      , and_dcpl_868 , and_dcpl_207 , and_dcpl_847});
  assign not_4418_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_46_nl = MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_re_0_14_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_39_16, {attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_3_39_16_mx0c1
      , and_dcpl_872 , and_dcpl_207 , and_dcpl_847});
  assign not_4417_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_47_nl = MUX1HOT_v_24_4_2(attention_2_1_16_16_4_4_k_proj_re_0_0_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16_mx0w1,
      attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_39_16, {attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_3_39_16_mx0c1
      , and_dcpl_876 , and_dcpl_207 , and_dcpl_847});
  assign not_4416_nl = ~ and_dcpl_619;
  assign GEMM_3D_FLOAT_LOOP_4_l_GEMM_3D_FLOAT_LOOP_4_l_mux_nl = MUX_s_1_2_2((z_out_5[1]),
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0]), APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c2);
  assign RMS_NORM_LOOP_2_2_mux_23_nl = MUX_s_1_16_2(1'b1, 1'b0, 1'b1, 1'b1, 1'b1,
      1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
      , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
  assign and_1810_nl = or_1907_cse & (fsm_output[4]);
  assign mux_2242_nl = MUX_s_1_2_2(nor_tmp_289, and_1810_nl, fsm_output[0]);
  assign mux_2243_nl = MUX_s_1_2_2((~ mux_2242_nl), nor_tmp_329, fsm_output[5]);
  assign mux_2244_nl = MUX_s_1_2_2((~ (fsm_output[5])), mux_2243_nl, fsm_output[3]);
  assign mux_2245_nl = MUX_s_1_2_2(mux_2244_nl, mux_tmp_1027, or_3039_cse);
  assign and_1254_nl = (~ mux_2245_nl) & and_dcpl_413;
  assign RMS_NORM_LOOP_1_1_mux1h_nl = MUX1HOT_s_1_3_2(RMS_NORM_LOOP_2_2_mux_23_nl,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1, (~ QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1),
      {and_dcpl_448 , and_1254_nl , and_dcpl_557});
  assign nor_1316_nl = ~((fsm_output[5]) | (or_1732_cse & (fsm_output[4:3]==2'b11)));
  assign and_1809_nl = (fsm_output[0]) & (fsm_output[1]) & (fsm_output[3]) & (fsm_output[4]);
  assign mux_2239_nl = MUX_s_1_2_2(nand_381_cse, and_1809_nl, fsm_output[5]);
  assign mux_2240_nl = MUX_s_1_2_2(nor_1316_nl, mux_2239_nl, fsm_output[2]);
  assign nor_1320_nl = ~((~ (fsm_output[8])) | (fsm_output[6]) | mux_2240_nl);
  assign or_3033_nl = (fsm_output[5:0]!=6'b101011);
  assign or_3032_nl = (fsm_output[5:0]!=6'b110100);
  assign mux_2238_nl = MUX_s_1_2_2(or_3033_nl, or_3032_nl, fsm_output[6]);
  assign nor_1321_nl = ~((fsm_output[8]) | mux_2238_nl);
  assign mux_2241_nl = MUX_s_1_2_2(nor_1320_nl, nor_1321_nl, fsm_output[7]);
  assign RMS_NORM_LOOP_1_1_or_nl = (RMS_NORM_LOOP_1_1_mux1h_nl & mux_2241_nl) | (and_dcpl_241
      & and_dcpl_293);
  assign GEMM_3D_FLOAT_LOOP_4_l_or_1_nl = and_dcpl_726 | APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c4;
  assign GEMM_3D_FLOAT_LOOP_4_l_mux1h_13_nl = MUX1HOT_s_1_3_2((z_out_5[0]), reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2,
      RMS_NORM_LOOP_1_1_or_nl, {GEMM_3D_FLOAT_LOOP_4_l_or_1_nl , APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c2
      , APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_mx0c3});
  assign and_939_nl = and_dcpl_732 & and_dcpl_875;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_26_nl = MUX1HOT_v_16_4_2(z_out_1,
      (rms_norm_16_div_cmp_z_oreg[15:0]), attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_2_0_0_sva_1_15_0, {and_939_nl , and_dcpl_876
      , and_dcpl_207 , and_dcpl_847});
  assign not_4471_nl = ~ and_dcpl_619;
  assign or_3191_nl = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b00) | (~ (fsm_output[0]))
      | mux_1639_cse;
  assign mux_1640_nl = MUX_s_1_2_2(or_2699_cse, or_3191_nl, and_1773_cse);
  assign or_3192_nl = (fsm_output[7]) | (~ mux_1640_nl);
  assign mux_1641_nl = MUX_s_1_2_2(nand_365_cse, or_3192_nl, fsm_output[6]);
  assign and_941_nl = and_dcpl_732 & and_dcpl_867;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_28_nl = MUX1HOT_v_16_4_2(z_out_1,
      (rms_norm_16_div_cmp_z_oreg[15:0]), attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_2_0_1_sva_1_15_0, {and_941_nl , and_dcpl_868
      , and_dcpl_207 , and_dcpl_847});
  assign not_4470_nl = ~ and_dcpl_619;
  assign or_3194_nl = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b01) | (~ (fsm_output[0]))
      | mux_1639_cse;
  assign mux_1643_nl = MUX_s_1_2_2(or_2699_cse, or_3194_nl, and_1773_cse);
  assign or_3195_nl = (fsm_output[7]) | (~ mux_1643_nl);
  assign mux_1644_nl = MUX_s_1_2_2(nand_365_cse, or_3195_nl, fsm_output[6]);
  assign and_958_nl = and_dcpl_732 & and_dcpl_879;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_40_nl = MUX1HOT_v_16_4_2(z_out_1,
      (rms_norm_16_div_cmp_z_oreg[15:0]), attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_3_0_3_sva_1_15_0, {and_958_nl , and_dcpl_880
      , and_dcpl_207 , and_dcpl_847});
  assign not_4464_nl = ~ and_dcpl_619;
  assign nand_81_nl = ~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2==2'b11) & (fsm_output[0])
      & (~ mux_1639_cse));
  assign mux_1726_nl = MUX_s_1_2_2(or_2699_cse, nand_81_nl, and_1773_cse);
  assign or_3197_nl = (fsm_output[7]) | (~ mux_1726_nl);
  assign mux_1727_nl = MUX_s_1_2_2(nand_365_cse, or_3197_nl, fsm_output[6]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_43_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_804);
  assign not_4458_nl = ~ and_dcpl_619;
  assign or_2491_nl = reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd!=3'b000);
  assign mux_1813_nl = MUX_s_1_2_2(mux_1812_cse, mux_806_cse, or_2491_nl);
  assign mux_1814_nl = MUX_s_1_2_2(or_2249_cse, mux_1813_nl, and_1773_cse);
  assign mux_1815_nl = MUX_s_1_2_2(mux_1814_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1816_nl = MUX_s_1_2_2(mux_1815_nl, or_1983_cse, fsm_output[5]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_42_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_796);
  assign not_4457_nl = ~ and_dcpl_619;
  assign or_2490_nl = (~ reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd!=3'b000);
  assign mux_1822_nl = MUX_s_1_2_2(mux_1812_cse, mux_806_cse, or_2490_nl);
  assign mux_1823_nl = MUX_s_1_2_2(or_2249_cse, mux_1822_nl, and_1773_cse);
  assign mux_1824_nl = MUX_s_1_2_2(mux_1823_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1825_nl = MUX_s_1_2_2(mux_1824_nl, or_1983_cse, fsm_output[5]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_41_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_776);
  assign not_4456_nl = ~ and_dcpl_619;
  assign nor_514_nl = ~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b10) | reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1
      | (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0])));
  assign mux_1831_nl = MUX_s_1_2_2(mux_806_cse, mux_1812_cse, nor_514_nl);
  assign mux_1832_nl = MUX_s_1_2_2(or_2249_cse, mux_1831_nl, and_1773_cse);
  assign mux_1833_nl = MUX_s_1_2_2(mux_1832_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1834_nl = MUX_s_1_2_2(mux_1833_nl, or_1983_cse, fsm_output[5]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_40_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_784);
  assign not_4455_nl = ~ and_dcpl_619;
  assign and_1727_nl = (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]==2'b10) & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1
      & (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]);
  assign mux_1840_nl = MUX_s_1_2_2(mux_806_cse, mux_1812_cse, and_1727_nl);
  assign mux_1841_nl = MUX_s_1_2_2(or_2249_cse, mux_1840_nl, and_1773_cse);
  assign mux_1842_nl = MUX_s_1_2_2(mux_1841_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1843_nl = MUX_s_1_2_2(mux_1842_nl, or_1983_cse, fsm_output[5]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_39_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_788);
  assign not_4454_nl = ~ and_dcpl_619;
  assign or_2653_nl = (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b11) | reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1
      | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]);
  assign mux_1849_nl = MUX_s_1_2_2(mux_1812_cse, mux_806_cse, or_2653_nl);
  assign mux_1850_nl = MUX_s_1_2_2(or_2249_cse, mux_1849_nl, and_1773_cse);
  assign mux_1851_nl = MUX_s_1_2_2(mux_1850_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1852_nl = MUX_s_1_2_2(mux_1851_nl, or_1983_cse, fsm_output[5]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_38_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_792);
  assign not_4453_nl = ~ and_dcpl_619;
  assign nand_369_nl = ~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]==2'b11) &
      reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 & (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0])));
  assign mux_1858_nl = MUX_s_1_2_2(mux_1812_cse, mux_806_cse, nand_369_nl);
  assign mux_1859_nl = MUX_s_1_2_2(or_2249_cse, mux_1858_nl, and_1773_cse);
  assign mux_1860_nl = MUX_s_1_2_2(mux_1859_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1861_nl = MUX_s_1_2_2(mux_1860_nl, or_1983_cse, fsm_output[5]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_37_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_800);
  assign not_4452_nl = ~ and_dcpl_619;
  assign and_1658_nl = (~ reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) & (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd==3'b111);
  assign mux_1867_nl = MUX_s_1_2_2(mux_806_cse, mux_1812_cse, and_1658_nl);
  assign mux_1868_nl = MUX_s_1_2_2(or_2249_cse, mux_1867_nl, and_1773_cse);
  assign mux_1869_nl = MUX_s_1_2_2(mux_1868_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1870_nl = MUX_s_1_2_2(mux_1869_nl, or_1983_cse, fsm_output[5]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_36_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_812);
  assign not_4451_nl = ~ and_dcpl_619;
  assign and_1733_nl = (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]==2'b11) & reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1
      & (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]) & (fsm_output[0]);
  assign mux_1874_nl = MUX_s_1_2_2(mux_806_cse, or_2249_cse, and_1733_nl);
  assign or_2664_nl = (~ (LINEAR_FORWARD_NO_MUL_LOOP_2_j_4_0_sva_1[4])) | (fsm_output[0]);
  assign mux_1873_nl = MUX_s_1_2_2(or_1983_cse, mux_806_cse, or_2664_nl);
  assign mux_1875_nl = MUX_s_1_2_2(mux_1874_nl, mux_1873_nl, fsm_output[1]);
  assign mux_1876_nl = MUX_s_1_2_2(or_2249_cse, mux_1875_nl, and_1773_cse);
  assign mux_1877_nl = MUX_s_1_2_2(mux_1876_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1878_nl = MUX_s_1_2_2(mux_1877_nl, or_1983_cse, fsm_output[5]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_35_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_959);
  assign not_4450_nl = ~ and_dcpl_619;
  assign nor_524_nl = ~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b00) | (~
      reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) | (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0])));
  assign mux_1884_nl = MUX_s_1_2_2(mux_806_cse, mux_1812_cse, nor_524_nl);
  assign mux_1885_nl = MUX_s_1_2_2(or_2249_cse, mux_1884_nl, and_1773_cse);
  assign mux_1886_nl = MUX_s_1_2_2(mux_1885_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1887_nl = MUX_s_1_2_2(mux_1886_nl, or_1983_cse, fsm_output[5]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_34_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_780);
  assign not_4449_nl = ~ and_dcpl_619;
  assign mux_1893_nl = MUX_s_1_2_2(mux_1812_cse, mux_806_cse, or_2671_cse);
  assign mux_1894_nl = MUX_s_1_2_2(or_2249_cse, mux_1893_nl, and_1773_cse);
  assign mux_1895_nl = MUX_s_1_2_2(mux_1894_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1896_nl = MUX_s_1_2_2(mux_1895_nl, or_1983_cse, fsm_output[5]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_33_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_772);
  assign not_4448_nl = ~ and_dcpl_619;
  assign or_2675_nl = (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b01) | (~
      reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]);
  assign mux_1902_nl = MUX_s_1_2_2(mux_1812_cse, mux_806_cse, or_2675_nl);
  assign mux_1903_nl = MUX_s_1_2_2(or_2249_cse, mux_1902_nl, and_1773_cse);
  assign mux_1904_nl = MUX_s_1_2_2(mux_1903_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1905_nl = MUX_s_1_2_2(mux_1904_nl, or_1983_cse, fsm_output[5]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_32_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_764);
  assign not_4447_nl = ~ and_dcpl_619;
  assign nor_441_nl = ~(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd!=3'b011));
  assign mux_1911_nl = MUX_s_1_2_2(mux_806_cse, mux_1812_cse, nor_441_nl);
  assign mux_1912_nl = MUX_s_1_2_2(or_2249_cse, mux_1911_nl, and_1773_cse);
  assign mux_1913_nl = MUX_s_1_2_2(mux_1912_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1914_nl = MUX_s_1_2_2(mux_1913_nl, or_1983_cse, fsm_output[5]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_31_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_754);
  assign not_4446_nl = ~ and_dcpl_619;
  assign and_1656_nl = reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 & (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd==3'b011);
  assign mux_1920_nl = MUX_s_1_2_2(mux_806_cse, mux_1812_cse, and_1656_nl);
  assign mux_1921_nl = MUX_s_1_2_2(or_2249_cse, mux_1920_nl, and_1773_cse);
  assign mux_1922_nl = MUX_s_1_2_2(mux_1921_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1923_nl = MUX_s_1_2_2(mux_1922_nl, or_1983_cse, fsm_output[5]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_30_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_760);
  assign not_4445_nl = ~ and_dcpl_619;
  assign mux_1929_nl = MUX_s_1_2_2(mux_1812_cse, mux_806_cse, or_2486_cse);
  assign mux_1930_nl = MUX_s_1_2_2(or_2249_cse, mux_1929_nl, and_1773_cse);
  assign mux_1931_nl = MUX_s_1_2_2(mux_1930_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1932_nl = MUX_s_1_2_2(mux_1931_nl, or_1983_cse, fsm_output[5]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux_29_nl = MUX_v_16_2_2(z_out, (rms_norm_16_div_cmp_z_oreg[15:0]),
      and_dcpl_768);
  assign not_4444_nl = ~ and_dcpl_619;
  assign or_2487_nl = (~ reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd!=3'b100);
  assign mux_1938_nl = MUX_s_1_2_2(mux_1812_cse, mux_806_cse, or_2487_nl);
  assign mux_1939_nl = MUX_s_1_2_2(or_2249_cse, mux_1938_nl, and_1773_cse);
  assign mux_1940_nl = MUX_s_1_2_2(mux_1939_nl, mux_1809_cse, fsm_output[4]);
  assign mux_1941_nl = MUX_s_1_2_2(mux_1940_nl, or_1983_cse, fsm_output[5]);
  assign and_1025_nl = and_dcpl_732 & and_dcpl_585 & and_dcpl_335;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_66_nl = MUX1HOT_v_16_4_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_v_proj_re_0_8_sva_2_15_0, attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0, {and_1025_nl , and_dcpl_983
      , and_dcpl_240 , and_dcpl_626});
  assign not_4563_nl = ~ and_dcpl_619;
  assign nor_533_nl = ~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 |
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1!=2'b00) | (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd));
  assign mux_1946_nl = MUX_s_1_2_2(mux_tmp_1945, mux_tmp_1943, nor_533_nl);
  assign and_1031_nl = and_dcpl_732 & and_dcpl_585 & and_dcpl_480;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_67_nl = MUX1HOT_v_16_4_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_v_proj_re_0_9_sva_2_15_0, attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0, {and_1031_nl , and_dcpl_983
      , and_dcpl_240 , and_dcpl_626});
  assign not_4564_nl = ~ and_dcpl_619;
  assign nor_535_nl = ~((~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2)
      | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1!=2'b00) | (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd));
  assign mux_1947_nl = MUX_s_1_2_2(mux_tmp_1945, mux_tmp_1943, nor_535_nl);
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_69_nl = MUX1HOT_v_8_7_2((drf_output_sdt_2_sva_15_0_mx0w0[15:8]),
      (attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_15_0[15:8]), (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0_mx0w1[15:8]),
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[15:8]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_15_8,
      (output_0_3_lpi_3_15_0[15:8]), (drf_output_sdt_3_sva_15_0_mx0w3[15:8]), {apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c1
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_626 , and_dcpl_207 , and_dcpl_739
      , apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c8});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_119_nl = MUX1HOT_v_8_7_2((drf_output_sdt_2_sva_15_0_mx0w0[7:0]),
      (attention_2_1_16_16_4_4_v_proj_re_0_3_sva_2_15_0[7:0]), (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0_mx0w1[7:0]),
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[7:0]), ({APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_7
      , APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_6
      , APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_5
      , APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_4
      , APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_3
      , APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_2
      , APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_1
      , APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_0}),
      (output_0_3_lpi_3_15_0[7:0]), (drf_output_sdt_3_sva_15_0_mx0w3[7:0]), {apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c1
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_626 , and_dcpl_207 , and_dcpl_739
      , apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0_mx0c8});
  assign not_4565_nl = ~ and_dcpl_619;
  assign nor_1203_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[7])) | (fsm_output[8]));
  assign nor_1204_nl = ~(and_1474_cse | (fsm_output[8:7]!=2'b01));
  assign mux_1970_nl = MUX_s_1_2_2(nor_1203_nl, nor_1204_nl, fsm_output[2]);
  assign nor_1201_nl = ~((~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd
      | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1 | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b11)))
      | (~ (fsm_output[0])) | (fsm_output[7]) | (~ (fsm_output[8])));
  assign nor_1202_nl = ~((fsm_output[8:7]!=2'b10));
  assign mux_1969_nl = MUX_s_1_2_2(nor_1201_nl, nor_1202_nl, fsm_output[1]);
  assign and_1749_nl = (fsm_output[2]) & mux_1969_nl;
  assign mux_1971_nl = MUX_s_1_2_2(mux_1970_nl, and_1749_nl, fsm_output[3]);
  assign and_1753_nl = (fsm_output[4]) & mux_1971_nl;
  assign nor_1206_nl = ~(((fsm_output[4:1]==4'b1111)) | (fsm_output[8:7]!=2'b10));
  assign mux_1972_nl = MUX_s_1_2_2(and_1753_nl, nor_1206_nl, fsm_output[5]);
  assign and_1754_nl = (fsm_output[3:2]==2'b11) & (~((~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd
      | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1]) | (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2)
      | (~ (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0])) | (fsm_output[1:0]!=2'b01)))
      | (fsm_output[8:7]!=2'b00)));
  assign mux_1967_nl = MUX_s_1_2_2(and_1754_nl, and_dcpl_26, fsm_output[4]);
  assign nor_1208_nl = ~((fsm_output[4]) | and_1638_cse | (fsm_output[8:7]!=2'b00));
  assign mux_1968_nl = MUX_s_1_2_2(mux_1967_nl, nor_1208_nl, fsm_output[5]);
  assign mux_1973_nl = MUX_s_1_2_2(mux_1972_nl, mux_1968_nl, fsm_output[6]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_70_nl = MUX1HOT_v_8_3_2((z_out[15:8]),
      (rms_norm_16_div_cmp_z_oreg[15:8]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm,
      {and_1042_ssc , and_dcpl_999 , and_dcpl_374});
  assign not_5074_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_128_nl = MUX1HOT_s_1_3_2((z_out[7]),
      (rms_norm_16_div_cmp_z_oreg[7]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm,
      {and_1042_ssc , and_dcpl_999 , and_dcpl_374});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_129_nl = MUX1HOT_s_1_3_2((z_out[6]),
      (rms_norm_16_div_cmp_z_oreg[6]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm,
      {and_1042_ssc , and_dcpl_999 , and_dcpl_374});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_130_nl = MUX1HOT_s_1_3_2((z_out[5]),
      (rms_norm_16_div_cmp_z_oreg[5]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm,
      {and_1042_ssc , and_dcpl_999 , and_dcpl_374});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_131_nl = MUX1HOT_s_1_3_2((z_out[4]),
      (rms_norm_16_div_cmp_z_oreg[4]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm,
      {and_1042_ssc , and_dcpl_999 , and_dcpl_374});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_132_nl = MUX1HOT_s_1_3_2((z_out[3]),
      (rms_norm_16_div_cmp_z_oreg[3]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm,
      {and_1042_ssc , and_dcpl_999 , and_dcpl_374});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_133_nl = MUX1HOT_s_1_3_2((z_out[2]),
      (rms_norm_16_div_cmp_z_oreg[2]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm,
      {and_1042_ssc , and_dcpl_999 , and_dcpl_374});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_134_nl = MUX1HOT_s_1_3_2((z_out[1]),
      (rms_norm_16_div_cmp_z_oreg[1]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm,
      {and_1042_ssc , and_dcpl_999 , and_dcpl_374});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_135_nl = MUX1HOT_s_1_3_2((z_out[0]),
      (rms_norm_16_div_cmp_z_oreg[0]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm,
      {and_1042_ssc , and_dcpl_999 , and_dcpl_374});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_71_nl = MUX1HOT_v_8_3_2((z_out_1[15:8]),
      (rms_norm_16_div_cmp_z_oreg[15:8]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_2_itm,
      {apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1 , and_dcpl_1003
      , and_dcpl_207});
  assign not_5066_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_120_nl = MUX1HOT_s_1_3_2((z_out_1[7]),
      (rms_norm_16_div_cmp_z_oreg[7]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_8_itm,
      {apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1 , and_dcpl_1003
      , and_dcpl_207});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_121_nl = MUX1HOT_s_1_3_2((z_out_1[6]),
      (rms_norm_16_div_cmp_z_oreg[6]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_9_itm,
      {apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1 , and_dcpl_1003
      , and_dcpl_207});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_122_nl = MUX1HOT_s_1_3_2((z_out_1[5]),
      (rms_norm_16_div_cmp_z_oreg[5]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_10_itm,
      {apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1 , and_dcpl_1003
      , and_dcpl_207});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_123_nl = MUX1HOT_s_1_3_2((z_out_1[4]),
      (rms_norm_16_div_cmp_z_oreg[4]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_11_itm,
      {apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1 , and_dcpl_1003
      , and_dcpl_207});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_124_nl = MUX1HOT_s_1_3_2((z_out_1[3]),
      (rms_norm_16_div_cmp_z_oreg[3]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_12_itm,
      {apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1 , and_dcpl_1003
      , and_dcpl_207});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_125_nl = MUX1HOT_s_1_3_2((z_out_1[2]),
      (rms_norm_16_div_cmp_z_oreg[2]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_13_itm,
      {apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1 , and_dcpl_1003
      , and_dcpl_207});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_126_nl = MUX1HOT_s_1_3_2((z_out_1[1]),
      (rms_norm_16_div_cmp_z_oreg[1]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_14_itm,
      {apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1 , and_dcpl_1003
      , and_dcpl_207});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_127_nl = MUX1HOT_s_1_3_2((z_out_1[0]),
      (rms_norm_16_div_cmp_z_oreg[0]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_APPLY_ROTARY_POS_EMB_LOOP_3_mux_15_itm,
      {apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_0_mx0c1 , and_dcpl_1003
      , and_dcpl_207});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_72_nl = MUX1HOT_v_16_5_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_v_proj_re_0_0_sva_2_15_0, z_out_1, output_0_0_lpi_3_15_0,
      drf_output_sdt_3_sva_15_0_mx0w3, {attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c1
      , and_dcpl_410 , and_dcpl_240 , and_dcpl_739 , attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0_mx0c6});
  assign not_4566_nl = ~ and_dcpl_619;
  assign mux_2010_nl = MUX_s_1_2_2(mux_304_cse, or_2457_cse, fsm_output[3]);
  assign nand_93_nl = ~((fsm_output[4]) & (~ mux_2010_nl));
  assign mux_2009_nl = MUX_s_1_2_2(mux_tmp_919, or_1197_cse, fsm_output[4]);
  assign mux_2011_nl = MUX_s_1_2_2(nand_93_nl, mux_2009_nl, fsm_output[5]);
  assign nand_92_nl = ~((fsm_output[3]) & (~((~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd
      | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1]) | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2
      | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0]) | (fsm_output[1:0]!=2'b01)))
      | (fsm_output[8:6]!=3'b001))));
  assign mux_2005_nl = MUX_s_1_2_2(mux_304_cse, or_2457_cse, and_1474_cse);
  assign and_1759_nl = or_3039_cse & (fsm_output[0]);
  assign mux_2002_nl = MUX_s_1_2_2(or_2457_cse, mux_tmp_919, and_1759_nl);
  assign mux_2003_nl = MUX_s_1_2_2(mux_2002_nl, mux_tmp_919, fsm_output[1]);
  assign mux_2006_nl = MUX_s_1_2_2(mux_2005_nl, mux_2003_nl, fsm_output[3]);
  assign mux_2007_nl = MUX_s_1_2_2(nand_92_nl, mux_2006_nl, fsm_output[4]);
  assign mux_2000_nl = MUX_s_1_2_2(mux_tmp_919, or_1197_cse, and_dcpl_65);
  assign or_2720_nl = and_dcpl_65 | (fsm_output[8:6]!=3'b100);
  assign mux_2001_nl = MUX_s_1_2_2(mux_2000_nl, or_2720_nl, fsm_output[4]);
  assign mux_2008_nl = MUX_s_1_2_2(mux_2007_nl, mux_2001_nl, fsm_output[5]);
  assign mux_2012_nl = MUX_s_1_2_2(mux_2011_nl, mux_2008_nl, fsm_output[2]);
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_73_nl = MUX1HOT_v_16_3_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_v_proj_re_0_7_sva_2_15_0, z_out, {attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0_mx0c1
      , and_dcpl_410 , and_dcpl_240});
  assign not_4567_nl = ~ and_dcpl_619;
  assign mux_2021_nl = MUX_s_1_2_2(mux_tmp_2015, mux_tmp_2013, fsm_output[3]);
  assign or_2733_nl = and_1762_cse | (fsm_output[7:6]!=2'b01);
  assign and_1763_nl = (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd) &
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1]) & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2
      & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0]) & (fsm_output[0]);
  assign mux_2018_nl = MUX_s_1_2_2(or_2733_nl, mux_tmp_2013, and_1763_nl);
  assign mux_2019_nl = MUX_s_1_2_2(mux_tmp_2015, mux_2018_nl, fsm_output[3]);
  assign mux_2016_nl = MUX_s_1_2_2(mux_tmp_2015, mux_tmp_2013, fsm_output[0]);
  assign mux_2017_nl = MUX_s_1_2_2(mux_2016_nl, or_tmp_914, fsm_output[3]);
  assign mux_2020_nl = MUX_s_1_2_2(mux_2019_nl, mux_2017_nl, fsm_output[1]);
  assign mux_2022_nl = MUX_s_1_2_2(mux_2021_nl, mux_2020_nl, fsm_output[2]);
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_nl = MUX_v_8_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[15:8]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[15:8]), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0[15:8]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0[15:8]), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3[15:8]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm[15:8]), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_15_8,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_15_8, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3[15:8]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm[15:8]), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_15_8,
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_8, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3[15:8]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm[15:8]), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_15_8,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_ftd, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_74_nl = MUX1HOT_v_8_9_2((drf_output_sdt_2_sva_15_0_mx0w0[15:8]),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_ftd, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_15_8,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_15_8, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_ftd, APPLY_ROTARY_POS_EMB_LOOP_6_mux_35_nl,
      output_0_1_lpi_3_15_8, (drf_output_sdt_3_sva_15_0_mx0w3[15:8]), {and_1055_ssc
      , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847
      , and_dcpl_583 , and_dcpl_739 , and_1059_ssc});
  assign not_5054_nl = ~ and_dcpl_619;
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_67_nl = MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[7]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[7]), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0[7]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0[7]), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3[7]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm[7]), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_7,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_7, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3[7]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm[7]), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_7,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3[7]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm[7]), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_7,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_117_nl = MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0[7]),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_7,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_7, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd, APPLY_ROTARY_POS_EMB_LOOP_6_mux_67_nl,
      output_0_1_lpi_3_7, (drf_output_sdt_3_sva_15_0_mx0w3[7]), {and_1055_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583
      , and_dcpl_739 , and_1059_ssc});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_88_nl = MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[6]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[6]), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0[6]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0[6]), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3[6]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm[6]), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_6,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_6, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3[6]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm[6]), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_6,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_1, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3[6]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm[6]), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_6,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_1, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_152_nl = MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0[6]),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_1, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_6,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_6, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_1, APPLY_ROTARY_POS_EMB_LOOP_6_mux_88_nl,
      output_0_1_lpi_3_6, (drf_output_sdt_3_sva_15_0_mx0w3[6]), {and_1055_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583
      , and_dcpl_739 , and_1059_ssc});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_89_nl = MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[5]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[5]), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0[5]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0[5]), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3[5]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm[5]), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_5,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_5, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3[5]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm[5]), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_5,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_2, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3[5]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm[5]), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_5,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_2, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_153_nl = MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0[5]),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_2, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_5,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_5, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_2, APPLY_ROTARY_POS_EMB_LOOP_6_mux_89_nl,
      output_0_1_lpi_3_5, (drf_output_sdt_3_sva_15_0_mx0w3[5]), {and_1055_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583
      , and_dcpl_739 , and_1059_ssc});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_90_nl = MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[4]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[4]), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0[4]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0[4]), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3[4]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm[4]), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_4,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_4, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3[4]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm[4]), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_4,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_3, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3[4]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm[4]), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_4,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_3, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_154_nl = MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0[4]),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_3, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_4,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_4, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_3, APPLY_ROTARY_POS_EMB_LOOP_6_mux_90_nl,
      output_0_1_lpi_3_4, (drf_output_sdt_3_sva_15_0_mx0w3[4]), {and_1055_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583
      , and_dcpl_739 , and_1059_ssc});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_91_nl = MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[3]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[3]), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0[3]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0[3]), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3[3]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm[3]), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_3,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_3, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3[3]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm[3]), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_3,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_4, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3[3]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm[3]), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_3,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_4, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_155_nl = MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0[3]),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_4, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_3,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_3, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_4, APPLY_ROTARY_POS_EMB_LOOP_6_mux_91_nl,
      output_0_1_lpi_3_3, (drf_output_sdt_3_sva_15_0_mx0w3[3]), {and_1055_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583
      , and_dcpl_739 , and_1059_ssc});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_92_nl = MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[2]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[2]), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0[2]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0[2]), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3[2]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm[2]), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_2,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_2, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3[2]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm[2]), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_2,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_5, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3[2]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm[2]), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_2,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_5, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_156_nl = MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0[2]),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_5, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_2,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_2, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_5, APPLY_ROTARY_POS_EMB_LOOP_6_mux_92_nl,
      output_0_1_lpi_3_2, (drf_output_sdt_3_sva_15_0_mx0w3[2]), {and_1055_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583
      , and_dcpl_739 , and_1059_ssc});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_93_nl = MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[1]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[1]), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0[1]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0[1]), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3[1]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm[1]), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_1,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_1, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3[1]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm[1]), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_1,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_6, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3[1]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm[1]), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_1,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_6, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_157_nl = MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0[1]),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_6, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_1,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_1, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_6, APPLY_ROTARY_POS_EMB_LOOP_6_mux_93_nl,
      output_0_1_lpi_3_1, (drf_output_sdt_3_sva_15_0_mx0w3[1]), {and_1055_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583
      , and_dcpl_739 , and_1059_ssc});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_94_nl = MUX_s_1_16_2((reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1[0]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[0]), (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0[0]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_15_0[0]), (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_0_lpi_3[0]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_1_0_1_lpi_3_dfm[0]), apply_rotary_pos_emb_1_4_4_rotated_k_1_0_2_1_lpi_3_0,
      apply_rotary_pos_emb_1_4_4_rotated_k_1_0_3_1_lpi_3_dfm_0, (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_0_lpi_3[0]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_2_0_1_lpi_3_dfm[0]), apply_rotary_pos_emb_1_4_4_rotated_k_2_0_2_1_lpi_3_0,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_15_0_1_ftd_7, (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_0_lpi_3[0]),
      (apply_rotary_pos_emb_1_4_4_rotated_k_3_0_1_lpi_3_dfm[0]), apply_rotary_pos_emb_1_4_4_rotated_k_3_0_2_1_lpi_3_0,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_7, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_158_nl = MUX1HOT_s_1_9_2((drf_output_sdt_2_sva_15_0_mx0w0[0]),
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_7, attention_2_1_16_16_4_4_v_proj_re_0_1_sva_2_0,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_mx0w1_0, apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0,
      reg_apply_rotary_pos_emb_1_4_4_rotated_k_3_0_3_1_lpi_3_dfm_15_0_1_ftd_7, APPLY_ROTARY_POS_EMB_LOOP_6_mux_94_nl,
      output_0_1_lpi_3_0, (drf_output_sdt_3_sva_15_0_mx0w3[0]), {and_1055_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583
      , and_dcpl_739 , and_1059_ssc});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_75_nl = MUX1HOT_v_3_6_2((drf_output_sdt_2_sva_15_0_mx0w0[15:13]),
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_13, attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_15_13,
      attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_15_13, apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_15_13,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_13, {and_1060_itm
      , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign not_4569_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_116_nl = MUX1HOT_v_5_7_2((drf_output_sdt_2_sva_15_0_mx0w0[12:8]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[12:8]), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0[12:8]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0[12:8]), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_12_8,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_12_8, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm[12:8]),
      {and_1060_itm , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207
      , and_dcpl_847 , and_dcpl_583});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_144_nl = MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0[7]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[7]), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0[7]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0[7]), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_7,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_7, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm[7]),
      {and_1060_itm , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207
      , and_dcpl_847 , and_dcpl_583});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_145_nl = MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0[6]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[6]), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0[6]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0[6]), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_6,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_6, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm[6]),
      {and_1060_itm , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207
      , and_dcpl_847 , and_dcpl_583});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_146_nl = MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0[5]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[5]), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0[5]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0[5]), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_5,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_5, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm[5]),
      {and_1060_itm , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207
      , and_dcpl_847 , and_dcpl_583});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_147_nl = MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0[4]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[4]), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0[4]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0[4]), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_4,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_4, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm[4]),
      {and_1060_itm , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207
      , and_dcpl_847 , and_dcpl_583});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_148_nl = MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0[3]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[3]), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0[3]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0[3]), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_3,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_3, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm[3]),
      {and_1060_itm , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207
      , and_dcpl_847 , and_dcpl_583});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_149_nl = MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0[2]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[2]), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0[2]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0[2]), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_2,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_2, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm[2]),
      {and_1060_itm , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207
      , and_dcpl_847 , and_dcpl_583});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_150_nl = MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0[1]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[1]), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0[1]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0[1]), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_1, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm[1]),
      {and_1060_itm , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207
      , and_dcpl_847 , and_dcpl_583});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_151_nl = MUX1HOT_s_1_7_2((drf_output_sdt_2_sva_15_0_mx0w0[0]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[0]), (attention_2_1_16_16_4_4_v_proj_re_0_10_sva_2_12_0[0]),
      (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_0_mx0w1_12_0[0]), apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_0_mx0w1_0,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_0, (APPLY_ROTARY_POS_EMB_LOOP_6_sinval_read_rom_sin_tab_rom_map_1_itm[0]),
      {and_1060_itm , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207
      , and_dcpl_847 , and_dcpl_583});
  assign not_5062_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_76_nl = MUX1HOT_v_8_6_2((drf_output_sdt_2_sva_15_0_mx0w0[15:8]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_8, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_15_8,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_15_8, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_15_8,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_8, {and_1062_ssc
      , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign not_5088_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_136_nl = MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0[7]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_7, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_7,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_7, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_7,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_7, {and_1062_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_137_nl = MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0[6]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_6, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_6,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_6, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_6,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_6, {and_1062_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_138_nl = MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0[5]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_5, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_5,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_5, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_5,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_5, {and_1062_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_139_nl = MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0[4]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_4, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_4,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_4, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_4,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_4, {and_1062_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_140_nl = MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0[3]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_3, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_3,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_3, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_3,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_3, {and_1062_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_141_nl = MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0[2]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_2, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_2,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_2, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_2,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_2, {and_1062_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_142_nl = MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0[1]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_1, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_1,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_1, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_1, {and_1062_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_143_nl = MUX1HOT_s_1_6_2((drf_output_sdt_2_sva_15_0_mx0w0[0]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_0, attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_0,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_0_mx0w1_0, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_0_mx0w1_0,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_0, {and_1062_ssc , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign and_1064_nl = and_dcpl_732 & and_dcpl_601;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_77_nl = MUX1HOT_v_16_6_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_v_proj_re_0_12_sva_2_15_0, attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0, attention_2_1_16_16_4_4_k_proj_2_0_0_lpi_3_15_0_mx0w6,
      attention_2_1_16_16_4_4_v_proj_0_0_0_sva_1_15_0, {and_1064_nl , and_dcpl_983
      , and_dcpl_240 , and_dcpl_626 , and_dcpl_207 , and_dcpl_213});
  assign not_4571_nl = ~ and_dcpl_619;
  assign nor_796_nl = ~((~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd)
      | (~ (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1])) | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2
      | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0]));
  assign mux_2038_nl = MUX_s_1_2_2(mux_tmp_1945, mux_tmp_1943, nor_796_nl);
  assign and_1066_nl = and_dcpl_732 & and_dcpl_595;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_78_nl = MUX1HOT_v_16_6_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_15_0,
      attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_0_0_1_sva_1_15_0, {and_1066_nl , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign not_4572_nl = ~ and_dcpl_619;
  assign and_1420_nl = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1])
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 & (~ (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0]));
  assign mux_2039_nl = MUX_s_1_2_2(mux_tmp_1945, mux_tmp_1943, and_1420_nl);
  assign and_1068_nl = and_dcpl_732 & and_dcpl_586;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_79_nl = MUX1HOT_v_16_6_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_re_0_14_sva_2_15_0,
      attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_0_0_2_sva_1_15_0, {and_1068_nl , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign not_4573_nl = ~ and_dcpl_619;
  assign and_1613_nl = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1])
      & (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2) & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0]);
  assign mux_2040_nl = MUX_s_1_2_2(mux_tmp_1945, mux_tmp_1943, and_1613_nl);
  assign and_1071_nl = and_dcpl_732 & and_dcpl_585 & and_dcpl_462;
  assign and_1074_nl = and_dcpl_743 & and_dcpl_740 & and_dcpl_854;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_80_nl = MUX1HOT_v_16_8_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_re_0_15_sva_2_15_0,
      attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_0_0_3_sva_1_15_0, output_0_15_lpi_3_15_0, drf_output_sdt_3_sva_15_0_mx0w3,
      {and_1071_nl , and_dcpl_1011 , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 ,
      and_dcpl_847 , and_dcpl_739 , and_1074_nl});
  assign not_4574_nl = ~ and_dcpl_619;
  assign or_2751_nl = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1])
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 & (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0]))
      | (~ (fsm_output[6])) | (fsm_output[8]);
  assign and_1660_nl = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2==2'b11)
      & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd & reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  assign mux_2045_nl = MUX_s_1_2_2(mux_tmp_121, or_tmp_464, and_1660_nl);
  assign mux_2046_nl = MUX_s_1_2_2(or_2751_nl, mux_2045_nl, fsm_output[4]);
  assign mux_2047_nl = MUX_s_1_2_2(or_tmp_464, mux_2046_nl, fsm_output[0]);
  assign mux_2048_nl = MUX_s_1_2_2(mux_2047_nl, mux_tmp_824, fsm_output[5]);
  assign mux_2049_nl = MUX_s_1_2_2(mux_2048_nl, mux_2025_cse, fsm_output[1]);
  assign mux_2051_nl = MUX_s_1_2_2(mux_2032_cse, mux_2049_nl, and_1773_cse);
  assign and_1075_nl = and_dcpl_732 & and_dcpl_598;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_81_nl = MUX1HOT_v_16_6_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_re_0_2_sva_2_15_0,
      attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0,
      attention_2_1_16_16_4_4_v_proj_1_0_0_sva_1_15_0_mx0w1, {and_1075_nl , attention_2_1_16_16_4_4_k_proj_re_or_cse
      , and_dcpl_983 , and_dcpl_240 , attention_2_1_16_16_4_4_k_proj_re_or_17_cse
      , and_dcpl_207});
  assign not_4575_nl = ~ and_dcpl_619;
  assign or_2753_nl = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1!=2'b01)
      | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd;
  assign mux_2052_nl = MUX_s_1_2_2(mux_tmp_1943, mux_tmp_1945, or_2753_nl);
  assign and_1081_nl = and_dcpl_732 & and_dcpl_610;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_82_nl = MUX1HOT_v_16_6_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_15_0,
      attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_1_0_1_sva_1_15_0, {and_1081_nl , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign not_4576_nl = ~ and_dcpl_619;
  assign or_2281_nl = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd | (~ (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1]))
      | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0]);
  assign mux_2053_nl = MUX_s_1_2_2(mux_tmp_1943, mux_tmp_1945, or_2281_nl);
  assign and_1083_nl = and_dcpl_732 & and_dcpl_616;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_83_nl = MUX1HOT_v_16_6_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_re_0_5_sva_2_15_0,
      attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_1_0_2_sva_1_15_0, {and_1083_nl , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign not_4577_nl = ~ and_dcpl_619;
  assign or_2292_nl = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd | (~ (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[1]))
      | (~ reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2) | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1[0]);
  assign mux_2054_nl = MUX_s_1_2_2(mux_tmp_1943, mux_tmp_1945, or_2292_nl);
  assign and_1086_nl = and_dcpl_732 & and_dcpl_591 & and_dcpl_486;
  assign attention_2_1_16_16_4_4_k_proj_re_mux1h_84_nl = MUX1HOT_v_16_6_2(drf_output_sdt_2_sva_15_0_mx0w0,
      attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0, attention_2_1_16_16_4_4_v_proj_re_0_6_sva_2_15_0,
      attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0_mx0w1, attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0_mx0w1,
      attention_2_1_16_16_4_4_v_proj_1_0_3_sva_1_15_0, {and_1086_nl , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847});
  assign not_4578_nl = ~ and_dcpl_619;
  assign or_2756_nl = reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_2 | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd_1!=2'b11)
      | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_2_j_4_0_sva_3_0_ftd;
  assign mux_2055_nl = MUX_s_1_2_2(mux_tmp_1943, mux_tmp_1945, or_2756_nl);
  assign or_2757_nl = (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b10)
      | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1;
  assign mux_2056_nl = MUX_s_1_2_2(nor_1026_cse, mux_tmp_1578, or_2757_nl);
  assign and_1089_nl = mux_2056_nl & (~ (fsm_output[8])) & and_dcpl_814;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_51_nl = MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_k_proj_re_0_2_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1,
      {and_1089_nl , and_dcpl_989 , and_dcpl_374});
  assign not_4414_nl = ~ and_dcpl_619;
  assign nor_1217_nl = ~((fsm_output[2]) | reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1
      | reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1 | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      | reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 | (~ (fsm_output[4])));
  assign mux_2057_nl = MUX_s_1_2_2(nor_1217_nl, and_1771_cse, fsm_output[1]);
  assign and_1090_nl = (fsm_output[0]) & mux_2057_nl;
  assign mux_2058_nl = MUX_s_1_2_2(and_1090_nl, (fsm_output[4]), fsm_output[3]);
  assign or_3200_nl = (fsm_output[7:6]!=2'b10) | mux_2058_nl;
  assign or_3201_nl = (~ (fsm_output[6])) | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_2059_nl = MUX_s_1_2_2(or_3200_nl, or_3201_nl, fsm_output[5]);
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_52_nl = MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_k_proj_re_0_3_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_k_proj_40_39_0_3_ctmp_sva_39_16_1,
      {apply_rotary_pos_emb_1_4_4_rotated_k_0_0_3_1_lpi_3_39_16_mx0c1 , and_dcpl_1003
      , and_dcpl_207});
  assign not_4413_nl = ~ and_dcpl_619;
  assign mux_2061_nl = MUX_s_1_2_2(and_dcpl_364, and_1771_cse, fsm_output[1]);
  assign or_2763_nl = (fsm_output[5]) | ((fsm_output[0]) & mux_2061_nl);
  assign mux_2062_nl = MUX_s_1_2_2(or_2763_nl, or_2699_cse, fsm_output[3]);
  assign or_2764_nl = (fsm_output[6]) | mux_2062_nl;
  assign mux_2063_nl = MUX_s_1_2_2(not_tmp_253, or_2764_nl, fsm_output[7]);
  assign or_2765_nl = reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd!=3'b001);
  assign mux_2064_nl = MUX_s_1_2_2(or_1983_cse, mux_tmp_1562, or_2765_nl);
  assign and_1097_nl = (~(mux_2064_nl | (fsm_output[8]))) & and_dcpl_748;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_53_nl = MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_q_proj_re_0_2_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1,
      {and_1097_nl , and_dcpl_999 , and_dcpl_374});
  assign not_4412_nl = ~ and_dcpl_619;
  assign nand_370_nl = ~((~((fsm_output[2:0]==3'b111))) & (fsm_output[4]));
  assign mux_2065_nl = MUX_s_1_2_2(nand_370_nl, or_tmp_330, fsm_output[3]);
  assign mux_2068_nl = MUX_s_1_2_2(mux_tmp_2067, mux_2065_nl, or_1880_cse);
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_54_nl = MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_q_proj_re_0_3_sva_1_39_16,
      (rms_norm_16_div_cmp_z_oreg[39:16]), APPLY_ROTARY_POS_EMB_LOOP_3_slc_attention_2_1_16_16_4_4_q_proj_40_39_0_2_ctmp_sva_39_16_1,
      {apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_39_16_mx0c1 , and_dcpl_959
      , and_dcpl_207});
  assign not_nl = ~ and_dcpl_619;
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_55_nl = MUX1HOT_v_24_3_2(attention_2_1_16_16_4_4_v_proj_re_0_4_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_4_sva_2_39_16, RESHAPE_2D_TO_3D_LOOP_3_1_slc_attention_2_1_16_16_4_4_k_proj_re_40_39_0_ctmp_sva_39_16_1,
      {and_dcpl_726 , and_dcpl_410 , and_dcpl_240});
  assign not_4579_nl = ~ and_dcpl_619;
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_36_nl = MUX_v_24_16_2(attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_39_16,
      attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_39_16, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_56_nl = MUX1HOT_v_24_9_2(attention_2_1_16_16_4_4_v_proj_re_0_13_sva_1_39_16,
      LINEAR_FORWARD_NO_MUL_LOOP_2_1_conc_1_mut_71_48_mx0w2, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_13_sva_2_39_16, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16_mx0w1,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16, apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_39_16_mx0w1,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_36_nl, LINEAR_FORWARD_NO_MUL_LOOP_2_3_conc_1_mut_71_48_mx0w3,
      {and_dcpl_726 , and_dcpl_257 , attention_2_1_16_16_4_4_k_proj_re_or_cse , and_dcpl_983
      , and_dcpl_240 , attention_2_1_16_16_4_4_k_proj_re_or_17_cse , and_dcpl_207
      , and_dcpl_583 , and_dcpl_265});
  assign not_4580_nl = ~ and_dcpl_619;
  assign LINEAR_FORWARD_NO_MUL_LOOP_2_mux_33_nl = MUX_v_24_16_2(attention_2_1_16_16_4_4_q_proj_re_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_1_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_re_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_3_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_re_0_4_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_5_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_re_0_6_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_7_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_re_0_8_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_9_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_re_0_10_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_11_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_re_0_12_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_13_sva_1_39_16, attention_2_1_16_16_4_4_q_proj_re_0_14_sva_1_39_16,
      attention_2_1_16_16_4_4_q_proj_re_0_15_sva_1_39_16, {reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd
      , reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_38_nl = MUX_v_24_16_2(attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_39_16,
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_39_16, attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_39_16, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign attention_2_1_16_16_4_4_v_proj_re_mux1h_57_nl = MUX1HOT_v_24_8_2(attention_2_1_16_16_4_4_v_proj_re_0_11_sva_1_39_16,
      LINEAR_FORWARD_NO_MUL_LOOP_2_mux_33_nl, attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16,
      attention_2_1_16_16_4_4_v_proj_re_0_11_sva_2_39_16, attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_39_16_mx0w1,
      apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16_mx0w1, apply_rotary_pos_emb_1_4_4_rotated_k_2_0_3_1_lpi_3_dfm_39_16,
      APPLY_ROTARY_POS_EMB_LOOP_6_mux_38_nl, {and_dcpl_726 , and_dcpl_257 , and_dcpl_1011
      , and_dcpl_983 , and_dcpl_240 , and_dcpl_207 , and_dcpl_847 , and_dcpl_583});
  assign not_4581_nl = ~ and_dcpl_619;
  assign QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_QUANTIZE_ACTIVATION_LOOP_3_nor_nl
      = ~((~ QUANTIZE_ACTIVATION_LOOP_3_quantized_value_clamped_acc_itm_25_1) | QUANTIZE_ACTIVATION_LOOP_3_nand_seb);
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_nl = MUX_v_8_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[15:8]),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1[15:8]), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_15_8,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_8, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3[15:8]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm[15:8]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_15_8, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3[15:8]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm[15:8]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd,
      ({apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_15_13 , apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_12_8}),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3[15:8]), (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm[15:8]),
      reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd, apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_15_8,
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_nl = MUX_v_8_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[15:8]),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_15_8, attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_8,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_ftd, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_15_8,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[15:8]), ({attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_15_13
      , (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[12:8])}), attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_15_8,
      (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[15:8]), (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[15:8]),
      (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0[15:8]), (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0[15:8]),
      (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[15:8]), (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[15:8]),
      (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0[15:8]), (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0[15:8]),
      {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_66_nl = MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[7]),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1[7]), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_7,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_7, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3[7]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm[7]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_7, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3[7]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm[7]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_7, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3[7]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm[7]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_7, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_74_nl = MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[6]),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1[6]), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_6,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_6, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3[6]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm[6]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_2,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_6, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3[6]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm[6]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_2,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_6, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3[6]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm[6]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_2,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_6, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_75_nl = MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[5]),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1[5]), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_5,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_5, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3[5]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm[5]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_3,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_5, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3[5]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm[5]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_3,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_5, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3[5]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm[5]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_3,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_5, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_76_nl = MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[4]),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1[4]), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_4,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_4, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3[4]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm[4]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_4,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_4, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3[4]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm[4]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_4,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_4, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3[4]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm[4]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_4,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_4, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_77_nl = MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[3]),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1[3]), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_3,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_3, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3[3]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm[3]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_5,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_3, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3[3]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm[3]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_5,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_3, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3[3]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm[3]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_5,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_3, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_78_nl = MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[2]),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1[2]), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_2,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_2, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3[2]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm[2]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_6,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_2, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3[2]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm[2]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_6,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_2, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3[2]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm[2]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_6,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_2, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_79_nl = MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[1]),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1[1]), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_1,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_1, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3[1]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm[1]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_7,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_1, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3[1]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm[1]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_7,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_1, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3[1]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm[1]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_7,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_1, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_80_nl = MUX_s_1_16_2((QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[0]),
      (reg_apply_rotary_pos_emb_1_4_4_rotated_q_0_0_1_ftd_1[0]), apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_0,
      apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_0, (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_0_lpi_3[0]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_1_0_1_lpi_3_dfm[0]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_1_0_2_1_lpi_3_15_0_ftd_8,
      apply_rotary_pos_emb_1_4_4_rotated_q_1_0_3_1_lpi_3_dfm_0, (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_0_lpi_3[0]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_2_0_1_lpi_3_dfm[0]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_2_1_lpi_3_15_0_ftd_8,
      apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_dfm_0, (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_0_lpi_3[0]),
      (apply_rotary_pos_emb_1_4_4_rotated_q_3_0_1_lpi_3_dfm[0]), reg_apply_rotary_pos_emb_1_4_4_rotated_q_3_0_2_1_lpi_3_15_0_ftd_8,
      apply_rotary_pos_emb_1_4_4_rotated_q_3_0_3_1_lpi_3_dfm_0, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_61_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[7]),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_7, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_7,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[7]), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[7]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_7, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[7]),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[7]), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0[7]),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0[7]), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[7]),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[7]), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0[7]),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0[7]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_81_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[6]),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_6, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_1,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_1, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_6,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[6]), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[6]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_6, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[6]),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[6]), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0[6]),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0[6]), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[6]),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[6]), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0[6]),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0[6]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_82_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[5]),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_5, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_2,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_2, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_5,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[5]), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[5]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_5, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[5]),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[5]), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0[5]),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0[5]), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[5]),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[5]), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0[5]),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0[5]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_83_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[4]),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_4, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_3,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_3, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_4,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[4]), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[4]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_4, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[4]),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[4]), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0[4]),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0[4]), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[4]),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[4]), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0[4]),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0[4]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_84_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[3]),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_3, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_4,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_4, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_3,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[3]), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[3]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_3, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[3]),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[3]), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0[3]),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0[3]), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[3]),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[3]), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0[3]),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0[3]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_85_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[2]),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_2, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_5,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_5, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_2,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[2]), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[2]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_2, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[2]),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[2]), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0[2]),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0[2]), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[2]),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[2]), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0[2]),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0[2]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_86_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[1]),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_1, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_6,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_6, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_1,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[1]), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[1]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_1, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[1]),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[1]), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0[1]),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0[1]), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[1]),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[1]), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0[1]),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0[1]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_87_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_k_proj_0_0_0_lpi_3_15_0[0]),
      attention_2_1_16_16_4_4_k_proj_0_0_1_sva_1_0, reg_attention_2_1_16_16_4_4_k_proj_0_0_2_sva_1_15_0_1_ftd_7,
      reg_attention_2_1_16_16_4_4_k_proj_0_0_3_sva_1_15_0_1_ftd_7, attention_2_1_16_16_4_4_k_proj_1_0_0_sva_1_0,
      (attention_2_1_16_16_4_4_k_proj_1_0_1_sva_1_15_0[0]), (attention_2_1_16_16_4_4_k_proj_1_0_2_sva_1_12_0[0]),
      attention_2_1_16_16_4_4_k_proj_1_0_3_sva_1_0, (attention_2_1_16_16_4_4_k_proj_2_0_0_sva_1_15_0[0]),
      (attention_2_1_16_16_4_4_k_proj_2_0_1_sva_1_15_0[0]), (attention_2_1_16_16_4_4_k_proj_2_0_2_sva_1_15_0[0]),
      (attention_2_1_16_16_4_4_k_proj_2_0_3_sva_1_15_0[0]), (attention_2_1_16_16_4_4_k_proj_3_0_0_sva_1_15_0[0]),
      (attention_2_1_16_16_4_4_k_proj_3_0_1_sva_1_15_0[0]), (attention_2_1_16_16_4_4_k_proj_3_0_2_sva_1_15_0[0]),
      (attention_2_1_16_16_4_4_k_proj_3_0_3_sva_1_15_0[0]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_32_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[15]),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[15]), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[15]),
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_15, (attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8[7]),
      (attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8[7]), (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8[7]),
      (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8[7]), (attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8[7]),
      (attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8[7]), (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8[7]),
      (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8[7]), (attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8[7]),
      (attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8[7]), (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8[7]),
      (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8[7]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_70_nl = MUX_v_3_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[14:12]),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[14:12]), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[14:12]),
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_14_12, (attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8[6:4]),
      (attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8[6:4]), (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8[6:4]),
      (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8[6:4]), (attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8[6:4]),
      (attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8[6:4]), (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8[6:4]),
      (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8[6:4]), (attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8[6:4]),
      (attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8[6:4]), (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8[6:4]),
      (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8[6:4]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_71_nl = MUX_v_3_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[11:9]),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[11:9]), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[11:9]),
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_11_9, (attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8[3:1]),
      (attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8[3:1]), (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8[3:1]),
      (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8[3:1]), (attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8[3:1]),
      (attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8[3:1]), (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8[3:1]),
      (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8[3:1]), (attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8[3:1]),
      (attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8[3:1]), (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8[3:1]),
      (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8[3:1]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_72_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[8]),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[8]), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[8]),
      attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_8, (attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_15_8[0]),
      (attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_15_8[0]), (attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_15_8[0]),
      (attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_15_8[0]), (attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_15_8[0]),
      (attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_15_8[0]), (attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_15_8[0]),
      (attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_15_8[0]), (attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_15_8[0]),
      (attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_15_8[0]), (attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_15_8[0]),
      (attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_15_8[0]), {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_50_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[7]),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[7]), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[7]),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[7]), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_7, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_7, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_7, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_7, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_7, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_7,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_7, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_51_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[6]),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[6]), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[6]),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[6]), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_6, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_6, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_6, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_6, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_6, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_6,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_6, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_52_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[5]),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[5]), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[5]),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[5]), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_5, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_5, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_5, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_5, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_5, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_5,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_5, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_53_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[4]),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[4]), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[4]),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[4]), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_4, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_4, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_4, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_4, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_4, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_4,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_4, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_54_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[3]),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[3]), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[3]),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[3]), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_3, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_3, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_3, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_3, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_3, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_3,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_3, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_55_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[2]),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[2]), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[2]),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[2]), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_2, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_2, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_2, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_2, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_2, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_2,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_2, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_56_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[1]),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[1]), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[1]),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[1]), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_1, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_1, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_1, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_1, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_1, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_1,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_1, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux_57_nl = MUX_s_1_16_2((attention_2_1_16_16_4_4_q_proj_0_0_0_lpi_3_15_0[0]),
      (attention_2_1_16_16_4_4_q_proj_0_0_1_sva_1_15_0[0]), (attention_2_1_16_16_4_4_q_proj_0_0_2_sva_1_15_0[0]),
      (attention_2_1_16_16_4_4_q_proj_0_0_3_sva_1_7_0[0]), attention_2_1_16_16_4_4_q_proj_1_0_0_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_1_0_1_sva_1_0, attention_2_1_16_16_4_4_q_proj_1_0_2_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_1_0_3_sva_1_0, attention_2_1_16_16_4_4_q_proj_2_0_0_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_2_0_1_sva_1_0, attention_2_1_16_16_4_4_q_proj_2_0_2_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_2_0_3_sva_1_0, attention_2_1_16_16_4_4_q_proj_3_0_0_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_3_0_1_sva_1_0, attention_2_1_16_16_4_4_q_proj_3_0_2_sva_1_0,
      attention_2_1_16_16_4_4_q_proj_3_0_3_sva_1_0, {reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1});
  assign APPLY_ROTARY_POS_EMB_LOOP_3_and_7_nl = (~ reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1)
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign APPLY_ROTARY_POS_EMB_LOOP_3_and_5_nl = reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1
      & reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1;
  assign mux_2129_nl = MUX_s_1_2_2((~ and_1570_cse), or_tmp_762, fsm_output[5]);
  assign mux_2130_nl = MUX_s_1_2_2(mux_2129_nl, or_tmp_682, fsm_output[3]);
  assign mux_2131_nl = MUX_s_1_2_2(and_1559_cse, (~ or_3137_cse), fsm_output[3]);
  assign attention_2_1_16_16_4_4_q_embed_or_nl = attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c1
      | (or_dcpl_996 & and_dcpl_204);
  assign attention_2_1_16_16_4_4_q_embed_and_33_nl = (~ or_dcpl_996) & and_dcpl_204;
  assign attention_2_1_16_16_4_4_q_embed_mux1h_40_nl = MUX1HOT_v_40_9_2(attention_2_1_16_16_4_4_q_embed_0_0_2_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1, APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_weights_3_0_0_sva_2, attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx1,
      attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx2, attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1,
      ({ATTN_2D_LOOP_3_mux_16_itm , ATTN_2D_LOOP_3_mux_17_itm}), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      {and_dcpl_346 , attention_2_1_16_16_4_4_q_embed_or_nl , attention_2_1_16_16_4_4_q_embed_and_33_nl
      , and_dcpl_348 , and_dcpl_349 , and_dcpl_351 , and_dcpl_1162 , and_dcpl_352
      , attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1_mx0c9});
  assign not_4510_nl = ~ mux_tmp_2153;
  assign attention_2_1_16_16_4_4_q_embed_mux1h_41_nl = MUX1HOT_v_40_6_2(attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1,
      attention_2_1_16_16_4_4_q_embed_0_0_3_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_weights_2_0_0_sva_2,
      attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx1, ({ATTN_2D_LOOP_3_mux_16_itm
      , ATTN_2D_LOOP_3_mux_17_itm}), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      {and_dcpl_346 , and_dcpl_204 , and_dcpl_348 , and_dcpl_351 , and_dcpl_352 ,
      attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1_mx0c7});
  assign not_4483_nl = ~ mux_tmp_2176;
  assign nor_1245_nl = ~((~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b00)
      | reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 | (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]))
      | (fsm_output[4:0]!=5'b10111))) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_2158_nl = MUX_s_1_2_2(mux_2157_cse, nor_1245_nl, fsm_output[5]);
  assign mux_2159_nl = MUX_s_1_2_2(nor_1239_cse, mux_2158_nl, fsm_output[7]);
  assign attention_2_1_16_16_4_4_q_embed_mux1h_42_nl = MUX1HOT_v_40_6_2(attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1,
      attention_2_1_16_16_4_4_q_embed_1_0_0_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_weights_3_0_1_sva_2,
      attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx1, ({ATTN_2D_LOOP_3_mux_16_itm
      , ATTN_2D_LOOP_3_mux_17_itm}), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      {and_dcpl_346 , and_dcpl_204 , and_dcpl_348 , and_dcpl_351 , and_dcpl_352 ,
      attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1_mx0c7});
  assign not_4482_nl = ~ mux_tmp_2176;
  assign nor_1256_nl = ~((~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b00)
      | (~ reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) | (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]))
      | (fsm_output[4:0]!=5'b10111))) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_2181_nl = MUX_s_1_2_2(mux_2157_cse, nor_1256_nl, fsm_output[5]);
  assign mux_2182_nl = MUX_s_1_2_2(nor_1239_cse, mux_2181_nl, fsm_output[7]);
  assign attention_2_1_16_16_4_4_q_embed_or_5_nl = attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c1
      | (or_dcpl_988 & and_dcpl_204);
  assign attention_2_1_16_16_4_4_q_embed_and_35_nl = (~ or_dcpl_988) & and_dcpl_204;
  assign attention_2_1_16_16_4_4_q_embed_mux1h_43_nl = MUX1HOT_v_40_9_2(attention_2_1_16_16_4_4_q_embed_1_0_1_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1, APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_1_sva_2, attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx1,
      attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx2, attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1,
      ({ATTN_2D_LOOP_3_mux_16_itm , ATTN_2D_LOOP_3_mux_17_itm}), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      {and_dcpl_346 , attention_2_1_16_16_4_4_q_embed_or_5_nl , attention_2_1_16_16_4_4_q_embed_and_35_nl
      , and_dcpl_348 , and_dcpl_349 , and_dcpl_351 , and_dcpl_1162 , and_dcpl_352
      , attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1_mx0c9});
  assign not_4511_nl = ~ mux_tmp_2153;
  assign attention_2_1_16_16_4_4_q_embed_mux1h_44_nl = MUX1HOT_v_40_6_2(attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1,
      attention_2_1_16_16_4_4_q_embed_1_0_2_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_weights_1_0_1_sva_2,
      attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx1, ({ATTN_2D_LOOP_3_mux_16_itm
      , ATTN_2D_LOOP_3_mux_17_itm}), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      {and_dcpl_346 , and_dcpl_204 , and_dcpl_348 , and_dcpl_351 , and_dcpl_352 ,
      attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1_mx0c7});
  assign not_4512_nl = ~ mux_tmp_2176;
  assign nor_1272_nl = ~((~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b01)
      | (~ reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0])
      | (fsm_output[4:0]!=5'b10111))) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_2197_nl = MUX_s_1_2_2(mux_2157_cse, nor_1272_nl, fsm_output[5]);
  assign mux_2198_nl = MUX_s_1_2_2(nor_1239_cse, mux_2197_nl, fsm_output[7]);
  assign attention_2_1_16_16_4_4_q_embed_mux1h_45_nl = MUX1HOT_v_40_6_2(attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1,
      attention_2_1_16_16_4_4_q_embed_1_0_3_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_weights_2_0_1_sva_2,
      attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx1, ({ATTN_2D_LOOP_3_mux_16_itm
      , ATTN_2D_LOOP_3_mux_17_itm}), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      {and_dcpl_346 , and_dcpl_204 , and_dcpl_348 , and_dcpl_351 , and_dcpl_352 ,
      attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1_mx0c7});
  assign not_4513_nl = ~ mux_tmp_2176;
  assign nor_1283_nl = ~((~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b01)
      | reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 | (~ (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]))
      | (fsm_output[4:0]!=5'b10111))) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_2203_nl = MUX_s_1_2_2(mux_2157_cse, nor_1283_nl, fsm_output[5]);
  assign mux_2204_nl = MUX_s_1_2_2(nor_1239_cse, mux_2203_nl, fsm_output[7]);
  assign attention_2_1_16_16_4_4_q_embed_mux1h_46_nl = MUX1HOT_v_40_6_2(attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1,
      attention_2_1_16_16_4_4_q_embed_2_0_0_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_weights_3_0_2_sva_2,
      attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx1, ({ATTN_2D_LOOP_3_mux_16_itm
      , ATTN_2D_LOOP_3_mux_17_itm}), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      {and_dcpl_346 , and_dcpl_204 , and_dcpl_348 , and_dcpl_351 , and_dcpl_352 ,
      attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1_mx0c7});
  assign not_4514_nl = ~ mux_tmp_2176;
  assign nor_1294_nl = ~(((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]==2'b01) &
      reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1 & (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0])
      & (fsm_output[4:0]==5'b10111)) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_2209_nl = MUX_s_1_2_2(mux_2157_cse, nor_1294_nl, fsm_output[5]);
  assign mux_2210_nl = MUX_s_1_2_2(nor_1239_cse, mux_2209_nl, fsm_output[7]);
  assign attention_2_1_16_16_4_4_q_embed_or_6_nl = attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c1
      | (or_dcpl_987 & and_dcpl_204);
  assign attention_2_1_16_16_4_4_q_embed_and_37_nl = (~ or_dcpl_987) & and_dcpl_204;
  assign attention_2_1_16_16_4_4_q_embed_mux1h_47_nl = MUX1HOT_v_40_9_2(attention_2_1_16_16_4_4_q_embed_2_0_1_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1, APPLY_ROTARY_POS_EMB_LOOP_6_acc_7_itm_55_16_1,
      attention_2_1_16_16_4_4_attn_weights_0_0_2_sva_2, attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx1,
      attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx2, attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1,
      ({ATTN_2D_LOOP_3_mux_16_itm , ATTN_2D_LOOP_3_mux_17_itm}), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      {and_dcpl_346 , attention_2_1_16_16_4_4_q_embed_or_6_nl , attention_2_1_16_16_4_4_q_embed_and_37_nl
      , and_dcpl_348 , and_dcpl_349 , and_dcpl_351 , and_dcpl_1162 , and_dcpl_352
      , attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1_mx0c9});
  assign not_4515_nl = ~ mux_tmp_2153;
  assign attention_2_1_16_16_4_4_q_embed_mux1h_48_nl = MUX1HOT_v_40_6_2(attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1,
      attention_2_1_16_16_4_4_q_embed_2_0_2_sva_1_mx0w1, attention_2_1_16_16_4_4_attn_weights_1_0_2_sva_2,
      attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx1, ({ATTN_2D_LOOP_3_mux_16_itm
      , ATTN_2D_LOOP_3_mux_17_itm}), RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_slc_71_32_1_ncse_sva,
      {and_dcpl_346 , and_dcpl_204 , and_dcpl_348 , and_dcpl_351 , and_dcpl_352 ,
      attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1_mx0c7});
  assign not_4516_nl = ~ mux_tmp_2176;
  assign nor_1310_nl = ~((~((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]!=2'b10)
      | (~ reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1) | (reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0])
      | (fsm_output[4:0]!=5'b10111))) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_2225_nl = MUX_s_1_2_2(mux_2157_cse, nor_1310_nl, fsm_output[5]);
  assign mux_2226_nl = MUX_s_1_2_2(nor_1239_cse, mux_2225_nl, fsm_output[7]);
  assign GEMM_3D_FLOAT_LOOP_3_not_28_nl = ~ GEMM_3D_FLOAT_LOOP_3_and_tmp_sva_mx0w0;
  assign GEMM_3D_FLOAT_LOOP_3_and_35_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1, GEMM_3D_FLOAT_LOOP_3_not_28_nl);
  assign GEMM_3D_FLOAT_LOOP_3_not_27_nl = ~ GEMM_3D_FLOAT_LOOP_3_and_tmp_11_sva_mx0w0;
  assign GEMM_3D_FLOAT_LOOP_3_and_34_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1, GEMM_3D_FLOAT_LOOP_3_not_27_nl);
  assign GEMM_3D_FLOAT_LOOP_3_not_26_nl = ~ GEMM_3D_FLOAT_LOOP_3_and_tmp_1_sva_mx0w0;
  assign GEMM_3D_FLOAT_LOOP_3_and_33_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1, GEMM_3D_FLOAT_LOOP_3_not_26_nl);
  assign GEMM_3D_FLOAT_LOOP_3_not_25_nl = ~ GEMM_3D_FLOAT_LOOP_3_and_tmp_10_sva_mx0w0;
  assign GEMM_3D_FLOAT_LOOP_3_and_32_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1, GEMM_3D_FLOAT_LOOP_3_not_25_nl);
  assign GEMM_3D_FLOAT_LOOP_3_not_24_nl = ~ GEMM_3D_FLOAT_LOOP_3_and_tmp_2_sva_mx0w0;
  assign GEMM_3D_FLOAT_LOOP_3_and_31_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1, GEMM_3D_FLOAT_LOOP_3_not_24_nl);
  assign GEMM_3D_FLOAT_LOOP_3_not_23_nl = ~ GEMM_3D_FLOAT_LOOP_3_and_tmp_9_sva_mx0w0;
  assign GEMM_3D_FLOAT_LOOP_3_and_30_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1, GEMM_3D_FLOAT_LOOP_3_not_23_nl);
  assign GEMM_3D_FLOAT_LOOP_3_not_22_nl = ~ GEMM_3D_FLOAT_LOOP_3_and_tmp_3_sva_mx0w0;
  assign GEMM_3D_FLOAT_LOOP_3_and_29_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1, GEMM_3D_FLOAT_LOOP_3_not_22_nl);
  assign GEMM_3D_FLOAT_LOOP_3_not_21_nl = ~ GEMM_3D_FLOAT_LOOP_3_and_tmp_8_sva_mx0w0;
  assign GEMM_3D_FLOAT_LOOP_3_and_28_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1, GEMM_3D_FLOAT_LOOP_3_not_21_nl);
  assign GEMM_3D_FLOAT_LOOP_3_not_20_nl = ~ GEMM_3D_FLOAT_LOOP_3_and_tmp_4_sva_mx0w2;
  assign GEMM_3D_FLOAT_LOOP_3_and_27_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1, GEMM_3D_FLOAT_LOOP_3_not_20_nl);
  assign GEMM_3D_FLOAT_LOOP_3_not_19_nl = ~ GEMM_3D_FLOAT_LOOP_3_and_tmp_7_sva_mx0w1;
  assign GEMM_3D_FLOAT_LOOP_3_and_26_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1, GEMM_3D_FLOAT_LOOP_3_not_19_nl);
  assign GEMM_3D_FLOAT_LOOP_3_not_18_nl = ~ GEMM_3D_FLOAT_LOOP_3_and_tmp_5_sva_mx0w2;
  assign GEMM_3D_FLOAT_LOOP_3_and_25_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1, GEMM_3D_FLOAT_LOOP_3_not_18_nl);
  assign GEMM_3D_FLOAT_LOOP_3_not_17_nl = ~ GEMM_3D_FLOAT_LOOP_3_and_tmp_6_sva_mx0w1;
  assign GEMM_3D_FLOAT_LOOP_3_and_24_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1, GEMM_3D_FLOAT_LOOP_3_not_17_nl);
  assign nor_1319_nl = ~((fsm_output[3]) | (fsm_output[5]) | or_tmp_1632);
  assign mux_2248_nl = MUX_s_1_2_2(mux_tmp_857, nor_1319_nl, fsm_output[6]);
  assign output_and_35_nl = or_dcpl_1155 & (~ and_dcpl_1232);
  assign output_and_39_nl = or_dcpl_1158 & (~ and_dcpl_1232);
  assign output_and_43_nl = or_dcpl_1160 & (~ and_dcpl_1232);
  assign output_and_47_nl = or_dcpl_1162 & (~ and_dcpl_1232);
  assign output_and_51_nl = or_dcpl_1165 & (~ and_dcpl_1232);
  assign output_and_55_nl = or_dcpl_1167 & (~ and_dcpl_1232);
  assign output_and_59_nl = or_dcpl_1169 & (~ and_dcpl_1232);
  assign output_and_63_nl = or_dcpl_1141 & (~ and_dcpl_1232);
  assign output_and_61_nl = or_dcpl_1170 & (~ and_dcpl_1232);
  assign output_and_57_nl = or_dcpl_1168 & (~ and_dcpl_1232);
  assign output_and_53_nl = or_dcpl_1166 & (~ and_dcpl_1232);
  assign output_and_49_nl = or_dcpl_1164 & (~ and_dcpl_1232);
  assign output_and_45_nl = or_dcpl_1161 & (~ and_dcpl_1232);
  assign output_and_41_nl = or_dcpl_1159 & (~ and_dcpl_1232);
  assign output_and_37_nl = or_dcpl_1156 & (~ and_dcpl_1232);
  assign output_and_33_nl = or_dcpl_1152 & (~ and_dcpl_1232);
  assign GEMM_3D_FLOAT_LOOP_4_l_mux1h_6_nl = MUX1HOT_s_1_3_2((z_out_3[1]), (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_k_2_0_sva_1[1]),
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[1]), {GEMM_3D_FLOAT_LOOP_4_l_or_2_cse
      , GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c3 , and_dcpl_193});
  assign operator_40_24_true_AC_TRN_AC_WRAP_or_nl = (acc_3_cse_40_1[3:0]!=4'b0000);
  assign nl_compute_sqrt_for_acc_3_nl = conv_u2s_3_4(z_out_12[3:1]) + 4'b1011;
  assign compute_sqrt_for_acc_3_nl = nl_compute_sqrt_for_acc_3_nl[3:0];
  assign RMS_NORM_LOOP_2_and_35_nl = RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_mux1h_itm &
      (~(RMS_NORM_LOOP_2_RMS_NORM_LOOP_2_nor_1_ssc_1 | RMS_NORM_LOOP_2_and_33_ssc_1));
  assign nor_658_nl = ~(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1 | reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1);
  assign RMS_NORM_LOOP_2_2_and_35_nl = RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_mux1h_itm
      & (~(RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_nor_1_ssc_1 | RMS_NORM_LOOP_2_2_and_33_ssc_1));
  assign mux_1258_nl = MUX_s_1_2_2(or_tmp_1664, mux_tmp_1245, and_1559_cse);
  assign mux_1254_nl = MUX_s_1_2_2(or_tmp_1066, mux_tmp_1237, fsm_output[5]);
  assign mux_1255_nl = MUX_s_1_2_2(mux_1254_nl, mux_tmp_1250, fsm_output[0]);
  assign mux_1256_nl = MUX_s_1_2_2(mux_tmp_1245, mux_1255_nl, fsm_output[2]);
  assign or_2167_nl = (fsm_output[8]) | mux_792_cse;
  assign mux_1252_nl = MUX_s_1_2_2(or_2167_nl, or_1197_cse, fsm_output[5]);
  assign mux_1247_nl = MUX_s_1_2_2(or_tmp_1066, or_1984_cse, fsm_output[5]);
  assign mux_1251_nl = MUX_s_1_2_2(mux_tmp_1250, mux_1247_nl, fsm_output[0]);
  assign mux_1253_nl = MUX_s_1_2_2(mux_1252_nl, mux_1251_nl, fsm_output[2]);
  assign mux_1257_nl = MUX_s_1_2_2(mux_1256_nl, mux_1253_nl, fsm_output[1]);
  assign mux_1259_nl = MUX_s_1_2_2(mux_1258_nl, mux_1257_nl, fsm_output[4]);
  assign or_3075_nl = (fsm_output[0]) | (fsm_output[2]);
  assign mux_1243_nl = MUX_s_1_2_2(mux_tmp_1240, mux_tmp_1238, or_3075_nl);
  assign nor_374_nl = ~(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd | reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      | (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2!=2'b00) | (~ (fsm_output[0])));
  assign mux_1241_nl = MUX_s_1_2_2(mux_tmp_1238, mux_tmp_1240, nor_374_nl);
  assign or_2162_nl = (fsm_output[5]) | mux_tmp_1237;
  assign mux_1239_nl = MUX_s_1_2_2(mux_tmp_1238, or_2162_nl, fsm_output[0]);
  assign mux_1242_nl = MUX_s_1_2_2(mux_1241_nl, mux_1239_nl, fsm_output[2]);
  assign mux_1244_nl = MUX_s_1_2_2(mux_1243_nl, mux_1242_nl, fsm_output[1]);
  assign mux_1246_nl = MUX_s_1_2_2(mux_tmp_1245, mux_1244_nl, fsm_output[4]);
  assign mux_1260_nl = MUX_s_1_2_2(mux_1259_nl, mux_1246_nl, fsm_output[3]);
  assign operator_40_24_true_AC_TRN_AC_WRAP_mux1h_nl = MUX1HOT_s_1_7_2(operator_40_24_true_AC_TRN_AC_WRAP_or_nl,
      (readslicef_4_1_3(compute_sqrt_for_acc_3_nl)), reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1,
      RMS_NORM_LOOP_2_and_35_nl, nor_658_nl, RMS_NORM_LOOP_2_2_and_35_nl, (~ QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_clamped_acc_itm_25_1),
      {rms_norm_16_variance_or_1_cse , and_dcpl_382 , (~ mux_1260_nl) , and_dcpl_344
      , and_dcpl_207 , and_dcpl_548 , and_dcpl_557});
  assign nor_1048_nl = ~((fsm_output[5]) | (fsm_output[0]) | (~ (fsm_output[4])));
  assign and_1603_nl = (fsm_output[5]) & (fsm_output[0]) & (fsm_output[1]) & (~ (fsm_output[4]));
  assign mux_1261_nl = MUX_s_1_2_2(nor_1048_nl, and_1603_nl, fsm_output[3]);
  assign QUANTIZE_ACTIVATION_LOOP_1_1_max_val_asn_GEMM_3D_FLOAT_LOOP_4_l_2_operator_40_24_true_AC_TRN_AC_WRAP_or_nl
      = (operator_40_24_true_AC_TRN_AC_WRAP_mux1h_nl & (~(mux_1261_nl & and_dcpl_390)))
      | and_dcpl_442;
  assign and_1256_nl = and_dcpl_191 & mux_tmp_787 & and_dcpl_293;
  assign mux_2246_nl = MUX_s_1_2_2(and_1762_cse, and_tmp_42, fsm_output[3]);
  assign nor_1318_nl = ~((fsm_output[3]) | (fsm_output[5]) | mux_tmp_1281);
  assign mux_2247_nl = MUX_s_1_2_2(mux_2246_nl, nor_1318_nl, fsm_output[6]);
  assign and_1257_nl = mux_2247_nl & GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c6;
  assign GEMM_3D_FLOAT_LOOP_4_l_mux1h_8_nl = MUX1HOT_s_1_7_2(QUANTIZE_ACTIVATION_LOOP_1_1_max_val_asn_GEMM_3D_FLOAT_LOOP_4_l_2_operator_40_24_true_AC_TRN_AC_WRAP_or_nl,
      (z_out_3[0]), (TRANSPOSE_LAST_TWO_DIMS_LOOP_3_k_2_0_sva_1[0]), (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]),
      CACHE_UPDATE_LOOP_2_1_acc_2_itm_2_1, reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1,
      CACHE_UPDATE_LOOP_2_acc_2_itm_2_1, {GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c0
      , GEMM_3D_FLOAT_LOOP_4_l_or_2_cse , GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_mx0c3
      , and_dcpl_193 , and_1256_nl , and_1257_nl , and_dcpl_316});
  assign CACHE_UPDATE_LOOP_3_mux1h_6_nl = MUX1HOT_s_1_3_2(reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0,
      reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd, (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[1]),
      {CACHE_UPDATE_LOOP_3_or_cse , CACHE_UPDATE_LOOP_3_or_1_cse , and_dcpl_1294});
  assign CACHE_UPDATE_LOOP_3_mux1h_7_nl = MUX1HOT_s_1_3_2(reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1,
      reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1, (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]),
      {CACHE_UPDATE_LOOP_3_or_cse , CACHE_UPDATE_LOOP_3_or_1_cse , and_dcpl_1294});
  assign nl_z_out_3 = conv_u2u_2_3({CACHE_UPDATE_LOOP_3_mux1h_6_nl , CACHE_UPDATE_LOOP_3_mux1h_7_nl})
      + 3'b001;
  assign z_out_3 = nl_z_out_3[2:0];
  assign nl_z_out_4 = conv_u2u_2_3({reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd
      , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1}) + 3'b001;
  assign z_out_4 = nl_z_out_4[2:0];
  assign GEMM_3D_FLOAT_LOOP_1_GEMM_3D_FLOAT_LOOP_1_mux_2_nl = MUX_s_1_2_2(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd, GEMM_3D_FLOAT_LOOP_1_or_ssc);
  assign GEMM_3D_FLOAT_LOOP_1_GEMM_3D_FLOAT_LOOP_1_mux_3_nl = MUX_s_1_2_2(reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1, GEMM_3D_FLOAT_LOOP_1_or_ssc);
  assign nl_z_out_5 = conv_u2u_2_3({GEMM_3D_FLOAT_LOOP_1_GEMM_3D_FLOAT_LOOP_1_mux_2_nl
      , GEMM_3D_FLOAT_LOOP_1_GEMM_3D_FLOAT_LOOP_1_mux_3_nl}) + 3'b001;
  assign z_out_5 = nl_z_out_5[2:0];
  assign nl_acc_3_cse_40_1 = ({reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd , reg_GEMM_3D_FLOAT_LOOP_4_1_mux_16_ftd_1})
      + ({reg_RMS_NORM_LOOP_1_1_slc_RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_mul_55_16_cse_1_slc
      , (APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm[39:16])});
  assign acc_3_cse_40_1 = nl_acc_3_cse_40_1[39:0];
  assign APPLY_ROTARY_POS_EMB_LOOP_6_APPLY_ROTARY_POS_EMB_LOOP_6_or_8_nl = (~(and_dcpl_1371
      | and_dcpl_1379)) | and_dcpl_1385;
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_36_nl = MUX1HOT_v_13_3_2(reg_apply_rotary_pos_emb_1_4_4_rotated_q_2_0_3_1_lpi_3_15_0_ftd_1,
      13'b0110100011101, 13'b1110001000111, {and_dcpl_1371 , and_dcpl_1379 , and_dcpl_1385});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_37_nl = MUX1HOT_v_24_3_2(for_for_strm_in_tmp_sva_25_2,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[39:16]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[39:16]),
      {and_dcpl_1371 , and_dcpl_1379 , and_dcpl_1385});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_38_nl = MUX1HOT_v_8_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[15:8]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[15:8]),
      {and_dcpl_1371 , and_dcpl_1379 , and_dcpl_1385});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_39_nl = MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_7,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[7]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[7]),
      {and_dcpl_1371 , and_dcpl_1379 , and_dcpl_1385});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_40_nl = MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_6,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[6]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[6]),
      {and_dcpl_1371 , and_dcpl_1379 , and_dcpl_1385});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_41_nl = MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_5,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[5]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[5]),
      {and_dcpl_1371 , and_dcpl_1379 , and_dcpl_1385});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_42_nl = MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_4,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[4]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[4]),
      {and_dcpl_1371 , and_dcpl_1379 , and_dcpl_1385});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_43_nl = MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_3,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[3]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[3]),
      {and_dcpl_1371 , and_dcpl_1379 , and_dcpl_1385});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_44_nl = MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_2,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[2]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[2]),
      {and_dcpl_1371 , and_dcpl_1379 , and_dcpl_1385});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_45_nl = MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_1,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[1]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[1]),
      {and_dcpl_1371 , and_dcpl_1379 , and_dcpl_1385});
  assign APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_46_nl = MUX1HOT_s_1_3_2(reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_33_itm_15_0_ftd_1_0,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[0]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[0]),
      {and_dcpl_1371 , and_dcpl_1379 , and_dcpl_1385});
  assign nl_z_out_9 = $signed(conv_u2s_20_21({(~ and_dcpl_1371) , 1'b0 , (~ and_dcpl_1371)
      , APPLY_ROTARY_POS_EMB_LOOP_6_APPLY_ROTARY_POS_EMB_LOOP_6_or_8_nl , (~ and_dcpl_1385)
      , (~ and_dcpl_1385) , (~ and_dcpl_1385) , APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_36_nl}))
      * $signed(({APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_37_nl , APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_38_nl
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_39_nl , APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_40_nl
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_41_nl , APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_42_nl
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_43_nl , APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_44_nl
      , APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_45_nl , APPLY_ROTARY_POS_EMB_LOOP_6_mux1h_46_nl}));
  assign z_out_9 = nl_z_out_9[59:0];
  assign RMS_NORM_LOOP_1_1_mux1h_134_nl = MUX1HOT_s_1_4_2((for_for_strm_in_tmp_sva_31_26[5]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[39]), QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39,
      (APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16[23]), {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_3_ssc
      , RMS_NORM_LOOP_1_1_or_1_ssc , and_dcpl_1415});
  assign RMS_NORM_LOOP_1_1_and_14_nl = RMS_NORM_LOOP_1_1_mux1h_134_nl & RMS_NORM_LOOP_1_1_nor_seb;
  assign RMS_NORM_LOOP_1_1_mux1h_135_nl = MUX1HOT_v_3_4_2((signext_3_1(for_for_strm_in_tmp_sva_31_26[5])),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[38:36]), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[38:36]),
      (APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16[22:20]), {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_3_ssc
      , RMS_NORM_LOOP_1_1_or_1_ssc , and_dcpl_1415});
  assign RMS_NORM_LOOP_1_1_and_15_nl = MUX_v_3_2_2(3'b000, RMS_NORM_LOOP_1_1_mux1h_135_nl,
      RMS_NORM_LOOP_1_1_nor_seb);
  assign RMS_NORM_LOOP_1_1_mux1h_136_nl = MUX1HOT_s_1_6_2((for_for_strm_in_tmp_sva_31_26[5]),
      attention_abs_qr_35_0_lpi_1_dfm_35, (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[35]),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[35]), (APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16[19]),
      attention_abs_4_qr_35_0_lpi_1_dfm_35, {and_dcpl_1393 , and_dcpl_1398 , RMS_NORM_LOOP_1_1_or_3_ssc
      , RMS_NORM_LOOP_1_1_or_1_ssc , and_dcpl_1415 , and_dcpl_1431});
  assign RMS_NORM_LOOP_1_1_mux1h_137_nl = MUX1HOT_v_6_6_2((signext_6_1(for_for_strm_in_tmp_sva_31_26[5])),
      (attention_abs_qr_35_0_lpi_1_dfm_34_0[34:29]), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[34:29]),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[34:29]), (APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16[18:13]),
      (attention_abs_4_qr_35_0_lpi_1_dfm_34_0[34:29]), {and_dcpl_1393 , and_dcpl_1398
      , RMS_NORM_LOOP_1_1_or_3_ssc , RMS_NORM_LOOP_1_1_or_1_ssc , and_dcpl_1415 ,
      and_dcpl_1431});
  assign RMS_NORM_LOOP_1_1_mux1h_138_nl = MUX1HOT_v_5_6_2((for_for_strm_in_tmp_sva_31_26[4:0]),
      (attention_abs_qr_35_0_lpi_1_dfm_34_0[28:24]), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[28:24]),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[28:24]), (APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16[12:8]),
      (attention_abs_4_qr_35_0_lpi_1_dfm_34_0[28:24]), {and_dcpl_1393 , and_dcpl_1398
      , RMS_NORM_LOOP_1_1_or_3_ssc , RMS_NORM_LOOP_1_1_or_1_ssc , and_dcpl_1415 ,
      and_dcpl_1431});
  assign RMS_NORM_LOOP_1_1_mux1h_139_nl = MUX1HOT_v_8_6_2((for_for_strm_in_tmp_sva_25_2[23:16]),
      (attention_abs_qr_35_0_lpi_1_dfm_34_0[23:16]), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[23:16]),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[23:16]), (APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_39_16[7:0]),
      (attention_abs_4_qr_35_0_lpi_1_dfm_34_0[23:16]), {and_dcpl_1393 , and_dcpl_1398
      , RMS_NORM_LOOP_1_1_or_3_ssc , RMS_NORM_LOOP_1_1_or_1_ssc , and_dcpl_1415 ,
      and_dcpl_1431});
  assign RMS_NORM_LOOP_1_1_mux1h_140_nl = MUX1HOT_v_8_6_2((for_for_strm_in_tmp_sva_25_2[15:8]),
      (attention_abs_qr_35_0_lpi_1_dfm_34_0[15:8]), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[15:8]),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[15:8]), reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd,
      (attention_abs_4_qr_35_0_lpi_1_dfm_34_0[15:8]), {and_dcpl_1393 , and_dcpl_1398
      , RMS_NORM_LOOP_1_1_or_3_ssc , RMS_NORM_LOOP_1_1_or_1_ssc , and_dcpl_1415 ,
      and_dcpl_1431});
  assign RMS_NORM_LOOP_1_1_mux1h_141_nl = MUX1HOT_v_8_6_2((for_for_strm_in_tmp_sva_25_2[7:0]),
      (attention_abs_qr_35_0_lpi_1_dfm_34_0[7:0]), (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[7:0]),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[7:0]), ({reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_7
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_6 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_5
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_4 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_3
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_2 , reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_1
      , reg_APPLY_ROTARY_POS_EMB_LOOP_6_mux_34_itm_15_0_ftd_1_0}), (attention_abs_4_qr_35_0_lpi_1_dfm_34_0[7:0]),
      {and_dcpl_1393 , and_dcpl_1398 , RMS_NORM_LOOP_1_1_or_3_ssc , RMS_NORM_LOOP_1_1_or_1_ssc
      , and_dcpl_1415 , and_dcpl_1431});
  assign RMS_NORM_LOOP_1_1_mux1h_142_nl = MUX1HOT_s_1_6_2((for_for_strm_in_tmp_sva_31_26[5]),
      (operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_17_16[1]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[39]), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd[2]),
      QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39, (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[39]),
      {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_4_itm , RMS_NORM_LOOP_1_1_or_2_ssc ,
      and_dcpl_1415 , and_dcpl_1420 , and_dcpl_1436});
  assign RMS_NORM_LOOP_1_1_and_16_nl = RMS_NORM_LOOP_1_1_mux1h_142_nl & (~ and_dcpl_1410)
      & (~ and_dcpl_1403);
  assign RMS_NORM_LOOP_1_1_mux1h_143_nl = MUX1HOT_v_15_6_2(({{9{for_for_strm_in_tmp_sva_31_26[5]}},
      for_for_strm_in_tmp_sva_31_26}), (signext_15_1(operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_17_16[1])),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[38:24]), (signext_15_1(reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd[2])),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[38:24]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[38:24]),
      {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_4_itm , RMS_NORM_LOOP_1_1_or_2_ssc ,
      and_dcpl_1415 , and_dcpl_1420 , and_dcpl_1436});
  assign RMS_NORM_LOOP_1_1_and_17_nl = RMS_NORM_LOOP_1_1_mux1h_143_nl & (signext_15_1(~
      and_dcpl_1410)) & (signext_15_1(~ and_dcpl_1403));
  assign RMS_NORM_LOOP_1_1_mux1h_144_nl = MUX1HOT_v_7_7_2((for_for_strm_in_tmp_sva_25_2[23:17]),
      (signext_7_1(operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_17_16[1])),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[23:17]), 7'b0000100, (signext_7_1(reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd[2])),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[23:17]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[23:17]),
      {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_4_itm , RMS_NORM_LOOP_1_1_or_2_ssc ,
      and_dcpl_1410 , and_dcpl_1415 , and_dcpl_1420 , and_dcpl_1436});
  assign not_5114_nl = ~ and_dcpl_1403;
  assign RMS_NORM_LOOP_1_1_and_18_nl = MUX_v_7_2_2(7'b0000000, RMS_NORM_LOOP_1_1_mux1h_144_nl,
      not_5114_nl);
  assign RMS_NORM_LOOP_1_1_mux1h_145_nl = MUX1HOT_s_1_6_2((for_for_strm_in_tmp_sva_25_2[16]),
      (operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_17_16[0]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[16]), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd[2]),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[16]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[16]),
      {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_4_itm , RMS_NORM_LOOP_1_1_or_2_ssc ,
      and_dcpl_1415 , and_dcpl_1420 , and_dcpl_1436});
  assign RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_3_nl = ~((~(RMS_NORM_LOOP_1_1_mux1h_145_nl
      | and_dcpl_1410)) | and_dcpl_1403);
  assign RMS_NORM_LOOP_1_1_mux1h_146_nl = MUX1HOT_s_1_6_2((for_for_strm_in_tmp_sva_25_2[15]),
      operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_itm_15,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[15]), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd[2]),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[15]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[15]),
      {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_4_itm , RMS_NORM_LOOP_1_1_or_2_ssc ,
      and_dcpl_1415 , and_dcpl_1420 , and_dcpl_1436});
  assign RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_4_nl = ~((~(RMS_NORM_LOOP_1_1_mux1h_146_nl
      | and_dcpl_1410)) | and_dcpl_1403);
  assign RMS_NORM_LOOP_1_1_mux1h_147_nl = MUX1HOT_v_2_6_2((for_for_strm_in_tmp_sva_25_2[14:13]),
      (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd[2:1]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[14:13]), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd[1:0]),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[14:13]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[14:13]),
      {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_4_itm , RMS_NORM_LOOP_1_1_or_2_ssc ,
      and_dcpl_1415 , and_dcpl_1420 , and_dcpl_1436});
  assign RMS_NORM_LOOP_1_1_and_19_nl = RMS_NORM_LOOP_1_1_mux1h_147_nl & (signext_2_1(~
      and_dcpl_1410)) & (signext_2_1(~ and_dcpl_1403));
  assign RMS_NORM_LOOP_1_1_mux1h_148_nl = MUX1HOT_s_1_6_2((for_for_strm_in_tmp_sva_25_2[12]),
      (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd[0]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[12]), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1[2]),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[12]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[12]),
      {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_4_itm , RMS_NORM_LOOP_1_1_or_2_ssc ,
      and_dcpl_1415 , and_dcpl_1420 , and_dcpl_1436});
  assign RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_5_nl = ~((~(RMS_NORM_LOOP_1_1_mux1h_148_nl
      | and_dcpl_1410)) | and_dcpl_1403);
  assign RMS_NORM_LOOP_1_1_mux1h_149_nl = MUX1HOT_v_2_7_2((for_for_strm_in_tmp_sva_25_2[11:10]),
      (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1[2:1]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[11:10]), 2'b01, (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1[1:0]),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[11:10]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[11:10]),
      {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_5_cse , RMS_NORM_LOOP_1_1_or_2_ssc ,
      and_dcpl_1410 , and_dcpl_1415 , and_dcpl_1420 , and_dcpl_1436});
  assign RMS_NORM_LOOP_1_1_mux1h_150_nl = MUX1HOT_s_1_6_2((for_for_strm_in_tmp_sva_25_2[9]),
      (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_1[0]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[9]), reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2,
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[9]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[9]),
      {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_5_cse , RMS_NORM_LOOP_1_1_or_2_ssc ,
      and_dcpl_1415 , and_dcpl_1420 , and_dcpl_1436});
  assign RMS_NORM_LOOP_1_1_and_20_nl = RMS_NORM_LOOP_1_1_mux1h_150_nl & (~ and_dcpl_1410);
  assign RMS_NORM_LOOP_1_1_mux1h_151_nl = MUX1HOT_s_1_6_2((for_for_strm_in_tmp_sva_25_2[8]),
      reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_2,
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[8]), (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3[7]),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[8]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[8]),
      {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_5_cse , RMS_NORM_LOOP_1_1_or_2_ssc ,
      and_dcpl_1415 , and_dcpl_1420 , and_dcpl_1436});
  assign RMS_NORM_LOOP_1_1_or_13_nl = RMS_NORM_LOOP_1_1_mux1h_151_nl | and_dcpl_1410;
  assign RMS_NORM_LOOP_1_1_mux1h_152_nl = MUX1HOT_v_2_7_2((for_for_strm_in_tmp_sva_25_2[7:6]),
      (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3[7:6]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[7:6]), 2'b01, (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3[6:5]),
      (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[7:6]), (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[7:6]),
      {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_5_cse , RMS_NORM_LOOP_1_1_or_2_ssc ,
      and_dcpl_1410 , and_dcpl_1415 , and_dcpl_1420 , and_dcpl_1436});
  assign RMS_NORM_LOOP_1_1_mux1h_153_nl = MUX1HOT_s_1_5_2((for_for_strm_in_tmp_sva_25_2[5]),
      (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3[5]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[5]), (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[5]),
      (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[5]), {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_5_cse
      , RMS_NORM_LOOP_1_1_or_2_ssc , and_dcpl_1420 , and_dcpl_1436});
  assign RMS_NORM_LOOP_1_1_or_14_nl = RMS_NORM_LOOP_1_1_mux1h_153_nl | and_dcpl_1415
      | and_dcpl_1410;
  assign RMS_NORM_LOOP_1_1_or_15_nl = and_dcpl_1398 | and_dcpl_1403 | and_dcpl_1415
      | and_dcpl_1431;
  assign RMS_NORM_LOOP_1_1_mux1h_154_nl = MUX1HOT_v_5_6_2((for_for_strm_in_tmp_sva_25_2[4:0]),
      (reg_operator_40_24_true_AC_TRN_AC_WRAP_1_slc_operator_40_24_true_AC_TRN_AC_WRAP_1_div_cmp_z_17_0_2_ftd_3[4:0]),
      (GEMM_3D_FLOAT_LOOP_4_1_mux_17_itm[4:0]), 5'b10001, (QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0[4:0]),
      (QUANTIZE_ACTIVATION_LOOP_1_1_scale_sva[4:0]), {and_dcpl_1393 , RMS_NORM_LOOP_1_1_or_15_nl
      , RMS_NORM_LOOP_1_1_or_2_ssc , and_dcpl_1410 , and_dcpl_1420 , and_dcpl_1436});
  assign nl_z_out_10 = $signed(({RMS_NORM_LOOP_1_1_and_14_nl , RMS_NORM_LOOP_1_1_and_15_nl
      , RMS_NORM_LOOP_1_1_mux1h_136_nl , RMS_NORM_LOOP_1_1_mux1h_137_nl , RMS_NORM_LOOP_1_1_mux1h_138_nl
      , RMS_NORM_LOOP_1_1_mux1h_139_nl , RMS_NORM_LOOP_1_1_mux1h_140_nl , RMS_NORM_LOOP_1_1_mux1h_141_nl}))
      * $signed(({RMS_NORM_LOOP_1_1_and_16_nl , RMS_NORM_LOOP_1_1_and_17_nl , RMS_NORM_LOOP_1_1_and_18_nl
      , RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_3_nl , RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_4_nl
      , RMS_NORM_LOOP_1_1_and_19_nl , RMS_NORM_LOOP_1_1_RMS_NORM_LOOP_1_1_nor_5_nl
      , RMS_NORM_LOOP_1_1_mux1h_149_nl , RMS_NORM_LOOP_1_1_and_20_nl , RMS_NORM_LOOP_1_1_or_13_nl
      , RMS_NORM_LOOP_1_1_mux1h_152_nl , RMS_NORM_LOOP_1_1_or_14_nl , RMS_NORM_LOOP_1_1_mux1h_154_nl}));
  assign z_out_10 = nl_z_out_10[63:0];
  assign TRANSPOSE_LAST_TWO_DIMS_LOOP_3_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_mux_2_nl =
      MUX_s_1_2_2(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd, reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd,
      and_dcpl_1447);
  assign TRANSPOSE_LAST_TWO_DIMS_LOOP_3_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_mux_3_nl =
      MUX_s_1_2_2(reg_GEMM_3D_FLOAT_LOOP_4_l_2_0_sva_1_0_ftd_1, reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1,
      and_dcpl_1447);
  assign nl_z_out_11 = conv_u2u_2_3({TRANSPOSE_LAST_TWO_DIMS_LOOP_3_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_mux_2_nl
      , TRANSPOSE_LAST_TWO_DIMS_LOOP_3_TRANSPOSE_LAST_TWO_DIMS_LOOP_3_mux_3_nl})
      + conv_u2u_2_3({reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1});
  assign z_out_11 = nl_z_out_11[2:0];
  assign nor_1397_nl = ~((fsm_output[2]) | (fsm_output[1]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1398_nl = ~((fsm_output[1]) | or_dcpl_959);
  assign and_2128_nl = (fsm_output[1]) & (fsm_output[4]) & (fsm_output[8]);
  assign mux_2303_nl = MUX_s_1_2_2(nor_1398_nl, and_2128_nl, fsm_output[2]);
  assign mux_2302_nl = MUX_s_1_2_2(nor_1397_nl, mux_2303_nl, fsm_output[3]);
  assign mux_2301_nl = MUX_s_1_2_2(mux_2302_nl, nor_1044_cse, fsm_output[6]);
  assign mux_2300_nl = MUX_s_1_2_2(mux_2301_nl, nor_1045_cse, fsm_output[7]);
  assign RMS_NORM_LOOP_2_2_or_1_nl = (and_dcpl_381 & (fsm_output[1:0]==2'b01) & and_dcpl_198)
      | (mux_2300_nl & (fsm_output[0]) & (~ (fsm_output[5])));
  assign RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_mux_1_nl = MUX_v_4_2_2(LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_1_3_0,
      ({reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2}), RMS_NORM_LOOP_2_2_or_1_nl);
  assign nl_z_out_12 = conv_u2u_4_5(RMS_NORM_LOOP_2_2_RMS_NORM_LOOP_2_2_mux_1_nl)
      + 5'b00001;
  assign z_out_12 = nl_z_out_12[4:0];
  assign and_2129_nl = (~ (fsm_output[8])) & (fsm_output[4]) & (fsm_output[1]) &
      (fsm_output[2]) & (fsm_output[0]) & (~ (fsm_output[3])) & (fsm_output[5]) &
      nor_973_cse;
  assign RMS_NORM_LOOP_2_2_mux_28_nl = MUX_v_53_2_2((APPLY_ROTARY_POS_EMB_LOOP_6_mul_3_itm[52:0]),
      (signext_53_52(APPLY_ROTARY_POS_EMB_LOOP_6_mul_2_itm[51:0])), and_2129_nl);
  assign nl_mul_3_nl = $signed(({QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_39
      , QUANTIZE_ACTIVATION_LOOP_3_1_quantized_value_mux_itm_38_0})) * $signed(RMS_NORM_LOOP_2_2_mux_28_nl);
  assign mul_3_nl = nl_mul_3_nl[71:0];
  assign z_out_13_71_28 = readslicef_72_44_28(mul_3_nl);
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_21_nl = MUX_v_2_2_2((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[2:1]),
      ({reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd , reg_APPLY_ROTARY_POS_EMB_LOOP_1_i_2_0_sva_1_0_ftd_1}),
      and_dcpl_1248);
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_22_nl = MUX_s_1_2_2((reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd[0]),
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd, and_dcpl_1248);
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_23_nl = MUX_s_1_2_2(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1,
      reg_GEMM_3D_FLOAT_LOOP_1_i_2_0_sva_1_0_ftd_1, and_dcpl_1248);
  assign z_out = MUX_v_16_16_2(attention_2_1_16_16_4_4_q_proj_re_0_0_lpi_4_15_0,
      attention_2_1_16_16_4_4_q_proj_re_0_1_lpi_4_15_0, ({apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_15_8
      , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_7 , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_6
      , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_5 , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_4
      , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_3 , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_2
      , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_1 , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_2_1_lpi_3_0}),
      attention_2_1_16_16_4_4_q_proj_re_0_3_lpi_4_15_0, attention_2_1_16_16_4_4_q_proj_re_0_4_lpi_4_15_0,
      attention_2_1_16_16_4_4_q_proj_re_0_5_lpi_4_15_0, attention_2_1_16_16_4_4_q_proj_re_0_6_lpi_4_15_0,
      attention_2_1_16_16_4_4_q_proj_re_0_7_lpi_4_15_0, attention_2_1_16_16_4_4_q_proj_re_0_8_lpi_4_15_0,
      attention_2_1_16_16_4_4_q_proj_re_0_9_lpi_4_15_0, attention_2_1_16_16_4_4_q_proj_re_0_10_lpi_4_15_0,
      attention_2_1_16_16_4_4_q_proj_re_0_11_lpi_4_15_0, attention_2_1_16_16_4_4_q_proj_re_0_12_lpi_4_15_0,
      attention_2_1_16_16_4_4_q_proj_re_0_13_lpi_4_15_0, attention_2_1_16_16_4_4_q_proj_re_0_14_lpi_4_15_0,
      attention_2_1_16_16_4_4_q_proj_re_0_15_lpi_4_15_0, {operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_21_nl
      , operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_22_nl , operator_40_24_true_AC_TRN_AC_WRAP_8_true_mux_23_nl});
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_22_nl = MUX_s_1_2_2(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd, and_dcpl_1261);
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_23_nl = MUX_s_1_2_2(reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1,
      reg_APPLY_ROTARY_POS_EMB_LOOP_6_k_2_0_sva_1_0_ftd_1, and_dcpl_1261);
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_24_nl = MUX_s_1_2_2((reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[1]),
      reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_0, and_dcpl_1261);
  assign operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_25_nl = MUX_s_1_2_2((reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]),
      reg_CACHE_UPDATE_LOOP_3_k_2_0_ftd_1, and_dcpl_1261);
  assign z_out_1 = MUX_v_16_16_2(attention_2_1_16_16_4_4_k_proj_re_0_0_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_1_lpi_4_15_0, apply_rotary_pos_emb_1_4_4_rotated_k_0_0_2_1_lpi_3_15_0,
      ({apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_15_8 , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_7
      , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_6 , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_5
      , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_4 , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_3
      , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_2 , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_1
      , apply_rotary_pos_emb_1_4_4_rotated_q_0_0_3_1_lpi_3_0}), attention_2_1_16_16_4_4_k_proj_re_0_4_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_5_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_6_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_7_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_8_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_9_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_10_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_11_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_12_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_13_lpi_4_15_0, attention_2_1_16_16_4_4_k_proj_re_0_14_lpi_4_15_0,
      attention_2_1_16_16_4_4_k_proj_re_0_15_lpi_4_15_0, {operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_22_nl
      , operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_23_nl , operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_24_nl
      , operator_40_24_true_AC_TRN_AC_WRAP_8_true_1_mux_25_nl});
  assign RMS_NORM_LOOP_2_2_mux_29_nl = MUX_v_3_2_2(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd,
      ({reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd , reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_1
      , (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[1])}), and_dcpl_1273);
  assign RMS_NORM_LOOP_2_2_mux_30_nl = MUX_s_1_2_2(reg_RMS_NORM_LOOP_2_2_i_4_0_sva_3_0_ftd_1,
      (reg_LINEAR_FORWARD_NO_MUL_LOOP_2_1_j_4_0_sva_3_0_ftd_2[0]), and_dcpl_1273);
  assign z_out_2 = MUX_v_40_16_2(attention_2_1_16_16_4_4_attn_output_2D_0_0_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_1_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_2_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_3_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_4_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_5_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_6_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_7_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_8_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_9_sva_1, attention_2_1_16_16_4_4_attn_output_2D_0_10_sva_1,
      attention_2_1_16_16_4_4_attn_output_2D_0_11_sva_1, attention_2_1_16_16_4_4_attn_output_3_0_0_lpi_3,
      attention_2_1_16_16_4_4_attn_output_3_0_1_lpi_3, attention_2_1_16_16_4_4_attn_output_3_0_2_lpi_3,
      attention_2_1_16_16_4_4_attn_output_3_0_3_lpi_3, {RMS_NORM_LOOP_2_2_mux_29_nl
      , RMS_NORM_LOOP_2_2_mux_30_nl});

  function automatic  MUX1HOT_s_1_13_2;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [12:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    MUX1HOT_s_1_13_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_5_2;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [4:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_6_2;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [5:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_7_2;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [6:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_8_2;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [7:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    MUX1HOT_s_1_8_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_9_2;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [8:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    MUX1HOT_s_1_9_2 = result;
  end
  endfunction


  function automatic [12:0] MUX1HOT_v_13_3_2;
    input [12:0] input_2;
    input [12:0] input_1;
    input [12:0] input_0;
    input [2:0] sel;
    reg [12:0] result;
  begin
    result = input_0 & {13{sel[0]}};
    result = result | (input_1 & {13{sel[1]}});
    result = result | (input_2 & {13{sel[2]}});
    MUX1HOT_v_13_3_2 = result;
  end
  endfunction


  function automatic [14:0] MUX1HOT_v_15_6_2;
    input [14:0] input_5;
    input [14:0] input_4;
    input [14:0] input_3;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [5:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | (input_1 & {15{sel[1]}});
    result = result | (input_2 & {15{sel[2]}});
    result = result | (input_3 & {15{sel[3]}});
    result = result | (input_4 & {15{sel[4]}});
    result = result | (input_5 & {15{sel[5]}});
    MUX1HOT_v_15_6_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_4_2;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [3:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    MUX1HOT_v_16_4_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_5_2;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [4:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    MUX1HOT_v_16_5_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_6_2;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [5:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    result = result | (input_5 & {16{sel[5]}});
    MUX1HOT_v_16_6_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_7_2;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [6:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    result = result | (input_5 & {16{sel[5]}});
    result = result | (input_6 & {16{sel[6]}});
    MUX1HOT_v_16_7_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_8_2;
    input [15:0] input_7;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [7:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    result = result | (input_5 & {16{sel[5]}});
    result = result | (input_6 & {16{sel[6]}});
    result = result | (input_7 & {16{sel[7]}});
    MUX1HOT_v_16_8_2 = result;
  end
  endfunction


  function automatic [20:0] MUX1HOT_v_21_5_2;
    input [20:0] input_4;
    input [20:0] input_3;
    input [20:0] input_2;
    input [20:0] input_1;
    input [20:0] input_0;
    input [4:0] sel;
    reg [20:0] result;
  begin
    result = input_0 & {21{sel[0]}};
    result = result | (input_1 & {21{sel[1]}});
    result = result | (input_2 & {21{sel[2]}});
    result = result | (input_3 & {21{sel[3]}});
    result = result | (input_4 & {21{sel[4]}});
    MUX1HOT_v_21_5_2 = result;
  end
  endfunction


  function automatic [21:0] MUX1HOT_v_22_5_2;
    input [21:0] input_4;
    input [21:0] input_3;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [4:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | (input_1 & {22{sel[1]}});
    result = result | (input_2 & {22{sel[2]}});
    result = result | (input_3 & {22{sel[3]}});
    result = result | (input_4 & {22{sel[4]}});
    MUX1HOT_v_22_5_2 = result;
  end
  endfunction


  function automatic [23:0] MUX1HOT_v_24_3_2;
    input [23:0] input_2;
    input [23:0] input_1;
    input [23:0] input_0;
    input [2:0] sel;
    reg [23:0] result;
  begin
    result = input_0 & {24{sel[0]}};
    result = result | (input_1 & {24{sel[1]}});
    result = result | (input_2 & {24{sel[2]}});
    MUX1HOT_v_24_3_2 = result;
  end
  endfunction


  function automatic [23:0] MUX1HOT_v_24_4_2;
    input [23:0] input_3;
    input [23:0] input_2;
    input [23:0] input_1;
    input [23:0] input_0;
    input [3:0] sel;
    reg [23:0] result;
  begin
    result = input_0 & {24{sel[0]}};
    result = result | (input_1 & {24{sel[1]}});
    result = result | (input_2 & {24{sel[2]}});
    result = result | (input_3 & {24{sel[3]}});
    MUX1HOT_v_24_4_2 = result;
  end
  endfunction


  function automatic [23:0] MUX1HOT_v_24_6_2;
    input [23:0] input_5;
    input [23:0] input_4;
    input [23:0] input_3;
    input [23:0] input_2;
    input [23:0] input_1;
    input [23:0] input_0;
    input [5:0] sel;
    reg [23:0] result;
  begin
    result = input_0 & {24{sel[0]}};
    result = result | (input_1 & {24{sel[1]}});
    result = result | (input_2 & {24{sel[2]}});
    result = result | (input_3 & {24{sel[3]}});
    result = result | (input_4 & {24{sel[4]}});
    result = result | (input_5 & {24{sel[5]}});
    MUX1HOT_v_24_6_2 = result;
  end
  endfunction


  function automatic [23:0] MUX1HOT_v_24_7_2;
    input [23:0] input_6;
    input [23:0] input_5;
    input [23:0] input_4;
    input [23:0] input_3;
    input [23:0] input_2;
    input [23:0] input_1;
    input [23:0] input_0;
    input [6:0] sel;
    reg [23:0] result;
  begin
    result = input_0 & {24{sel[0]}};
    result = result | (input_1 & {24{sel[1]}});
    result = result | (input_2 & {24{sel[2]}});
    result = result | (input_3 & {24{sel[3]}});
    result = result | (input_4 & {24{sel[4]}});
    result = result | (input_5 & {24{sel[5]}});
    result = result | (input_6 & {24{sel[6]}});
    MUX1HOT_v_24_7_2 = result;
  end
  endfunction


  function automatic [23:0] MUX1HOT_v_24_8_2;
    input [23:0] input_7;
    input [23:0] input_6;
    input [23:0] input_5;
    input [23:0] input_4;
    input [23:0] input_3;
    input [23:0] input_2;
    input [23:0] input_1;
    input [23:0] input_0;
    input [7:0] sel;
    reg [23:0] result;
  begin
    result = input_0 & {24{sel[0]}};
    result = result | (input_1 & {24{sel[1]}});
    result = result | (input_2 & {24{sel[2]}});
    result = result | (input_3 & {24{sel[3]}});
    result = result | (input_4 & {24{sel[4]}});
    result = result | (input_5 & {24{sel[5]}});
    result = result | (input_6 & {24{sel[6]}});
    result = result | (input_7 & {24{sel[7]}});
    MUX1HOT_v_24_8_2 = result;
  end
  endfunction


  function automatic [23:0] MUX1HOT_v_24_9_2;
    input [23:0] input_8;
    input [23:0] input_7;
    input [23:0] input_6;
    input [23:0] input_5;
    input [23:0] input_4;
    input [23:0] input_3;
    input [23:0] input_2;
    input [23:0] input_1;
    input [23:0] input_0;
    input [8:0] sel;
    reg [23:0] result;
  begin
    result = input_0 & {24{sel[0]}};
    result = result | (input_1 & {24{sel[1]}});
    result = result | (input_2 & {24{sel[2]}});
    result = result | (input_3 & {24{sel[3]}});
    result = result | (input_4 & {24{sel[4]}});
    result = result | (input_5 & {24{sel[5]}});
    result = result | (input_6 & {24{sel[6]}});
    result = result | (input_7 & {24{sel[7]}});
    result = result | (input_8 & {24{sel[8]}});
    MUX1HOT_v_24_9_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_6_2;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [5:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    MUX1HOT_v_2_6_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_7_2;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [6:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    MUX1HOT_v_2_7_2 = result;
  end
  endfunction


  function automatic [33:0] MUX1HOT_v_34_7_2;
    input [33:0] input_6;
    input [33:0] input_5;
    input [33:0] input_4;
    input [33:0] input_3;
    input [33:0] input_2;
    input [33:0] input_1;
    input [33:0] input_0;
    input [6:0] sel;
    reg [33:0] result;
  begin
    result = input_0 & {34{sel[0]}};
    result = result | (input_1 & {34{sel[1]}});
    result = result | (input_2 & {34{sel[2]}});
    result = result | (input_3 & {34{sel[3]}});
    result = result | (input_4 & {34{sel[4]}});
    result = result | (input_5 & {34{sel[5]}});
    result = result | (input_6 & {34{sel[6]}});
    MUX1HOT_v_34_7_2 = result;
  end
  endfunction


  function automatic [37:0] MUX1HOT_v_38_5_2;
    input [37:0] input_4;
    input [37:0] input_3;
    input [37:0] input_2;
    input [37:0] input_1;
    input [37:0] input_0;
    input [4:0] sel;
    reg [37:0] result;
  begin
    result = input_0 & {38{sel[0]}};
    result = result | (input_1 & {38{sel[1]}});
    result = result | (input_2 & {38{sel[2]}});
    result = result | (input_3 & {38{sel[3]}});
    result = result | (input_4 & {38{sel[4]}});
    MUX1HOT_v_38_5_2 = result;
  end
  endfunction


  function automatic [38:0] MUX1HOT_v_39_10_2;
    input [38:0] input_9;
    input [38:0] input_8;
    input [38:0] input_7;
    input [38:0] input_6;
    input [38:0] input_5;
    input [38:0] input_4;
    input [38:0] input_3;
    input [38:0] input_2;
    input [38:0] input_1;
    input [38:0] input_0;
    input [9:0] sel;
    reg [38:0] result;
  begin
    result = input_0 & {39{sel[0]}};
    result = result | (input_1 & {39{sel[1]}});
    result = result | (input_2 & {39{sel[2]}});
    result = result | (input_3 & {39{sel[3]}});
    result = result | (input_4 & {39{sel[4]}});
    result = result | (input_5 & {39{sel[5]}});
    result = result | (input_6 & {39{sel[6]}});
    result = result | (input_7 & {39{sel[7]}});
    result = result | (input_8 & {39{sel[8]}});
    result = result | (input_9 & {39{sel[9]}});
    MUX1HOT_v_39_10_2 = result;
  end
  endfunction


  function automatic [38:0] MUX1HOT_v_39_13_2;
    input [38:0] input_12;
    input [38:0] input_11;
    input [38:0] input_10;
    input [38:0] input_9;
    input [38:0] input_8;
    input [38:0] input_7;
    input [38:0] input_6;
    input [38:0] input_5;
    input [38:0] input_4;
    input [38:0] input_3;
    input [38:0] input_2;
    input [38:0] input_1;
    input [38:0] input_0;
    input [12:0] sel;
    reg [38:0] result;
  begin
    result = input_0 & {39{sel[0]}};
    result = result | (input_1 & {39{sel[1]}});
    result = result | (input_2 & {39{sel[2]}});
    result = result | (input_3 & {39{sel[3]}});
    result = result | (input_4 & {39{sel[4]}});
    result = result | (input_5 & {39{sel[5]}});
    result = result | (input_6 & {39{sel[6]}});
    result = result | (input_7 & {39{sel[7]}});
    result = result | (input_8 & {39{sel[8]}});
    result = result | (input_9 & {39{sel[9]}});
    result = result | (input_10 & {39{sel[10]}});
    result = result | (input_11 & {39{sel[11]}});
    result = result | (input_12 & {39{sel[12]}});
    MUX1HOT_v_39_13_2 = result;
  end
  endfunction


  function automatic [38:0] MUX1HOT_v_39_3_2;
    input [38:0] input_2;
    input [38:0] input_1;
    input [38:0] input_0;
    input [2:0] sel;
    reg [38:0] result;
  begin
    result = input_0 & {39{sel[0]}};
    result = result | (input_1 & {39{sel[1]}});
    result = result | (input_2 & {39{sel[2]}});
    MUX1HOT_v_39_3_2 = result;
  end
  endfunction


  function automatic [38:0] MUX1HOT_v_39_5_2;
    input [38:0] input_4;
    input [38:0] input_3;
    input [38:0] input_2;
    input [38:0] input_1;
    input [38:0] input_0;
    input [4:0] sel;
    reg [38:0] result;
  begin
    result = input_0 & {39{sel[0]}};
    result = result | (input_1 & {39{sel[1]}});
    result = result | (input_2 & {39{sel[2]}});
    result = result | (input_3 & {39{sel[3]}});
    result = result | (input_4 & {39{sel[4]}});
    MUX1HOT_v_39_5_2 = result;
  end
  endfunction


  function automatic [38:0] MUX1HOT_v_39_8_2;
    input [38:0] input_7;
    input [38:0] input_6;
    input [38:0] input_5;
    input [38:0] input_4;
    input [38:0] input_3;
    input [38:0] input_2;
    input [38:0] input_1;
    input [38:0] input_0;
    input [7:0] sel;
    reg [38:0] result;
  begin
    result = input_0 & {39{sel[0]}};
    result = result | (input_1 & {39{sel[1]}});
    result = result | (input_2 & {39{sel[2]}});
    result = result | (input_3 & {39{sel[3]}});
    result = result | (input_4 & {39{sel[4]}});
    result = result | (input_5 & {39{sel[5]}});
    result = result | (input_6 & {39{sel[6]}});
    result = result | (input_7 & {39{sel[7]}});
    MUX1HOT_v_39_8_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_5_2;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [4:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    MUX1HOT_v_3_5_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_6_2;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [5:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    result = result | (input_5 & {3{sel[5]}});
    MUX1HOT_v_3_6_2 = result;
  end
  endfunction


  function automatic [39:0] MUX1HOT_v_40_10_2;
    input [39:0] input_9;
    input [39:0] input_8;
    input [39:0] input_7;
    input [39:0] input_6;
    input [39:0] input_5;
    input [39:0] input_4;
    input [39:0] input_3;
    input [39:0] input_2;
    input [39:0] input_1;
    input [39:0] input_0;
    input [9:0] sel;
    reg [39:0] result;
  begin
    result = input_0 & {40{sel[0]}};
    result = result | (input_1 & {40{sel[1]}});
    result = result | (input_2 & {40{sel[2]}});
    result = result | (input_3 & {40{sel[3]}});
    result = result | (input_4 & {40{sel[4]}});
    result = result | (input_5 & {40{sel[5]}});
    result = result | (input_6 & {40{sel[6]}});
    result = result | (input_7 & {40{sel[7]}});
    result = result | (input_8 & {40{sel[8]}});
    result = result | (input_9 & {40{sel[9]}});
    MUX1HOT_v_40_10_2 = result;
  end
  endfunction


  function automatic [39:0] MUX1HOT_v_40_11_2;
    input [39:0] input_10;
    input [39:0] input_9;
    input [39:0] input_8;
    input [39:0] input_7;
    input [39:0] input_6;
    input [39:0] input_5;
    input [39:0] input_4;
    input [39:0] input_3;
    input [39:0] input_2;
    input [39:0] input_1;
    input [39:0] input_0;
    input [10:0] sel;
    reg [39:0] result;
  begin
    result = input_0 & {40{sel[0]}};
    result = result | (input_1 & {40{sel[1]}});
    result = result | (input_2 & {40{sel[2]}});
    result = result | (input_3 & {40{sel[3]}});
    result = result | (input_4 & {40{sel[4]}});
    result = result | (input_5 & {40{sel[5]}});
    result = result | (input_6 & {40{sel[6]}});
    result = result | (input_7 & {40{sel[7]}});
    result = result | (input_8 & {40{sel[8]}});
    result = result | (input_9 & {40{sel[9]}});
    result = result | (input_10 & {40{sel[10]}});
    MUX1HOT_v_40_11_2 = result;
  end
  endfunction


  function automatic [39:0] MUX1HOT_v_40_3_2;
    input [39:0] input_2;
    input [39:0] input_1;
    input [39:0] input_0;
    input [2:0] sel;
    reg [39:0] result;
  begin
    result = input_0 & {40{sel[0]}};
    result = result | (input_1 & {40{sel[1]}});
    result = result | (input_2 & {40{sel[2]}});
    MUX1HOT_v_40_3_2 = result;
  end
  endfunction


  function automatic [39:0] MUX1HOT_v_40_6_2;
    input [39:0] input_5;
    input [39:0] input_4;
    input [39:0] input_3;
    input [39:0] input_2;
    input [39:0] input_1;
    input [39:0] input_0;
    input [5:0] sel;
    reg [39:0] result;
  begin
    result = input_0 & {40{sel[0]}};
    result = result | (input_1 & {40{sel[1]}});
    result = result | (input_2 & {40{sel[2]}});
    result = result | (input_3 & {40{sel[3]}});
    result = result | (input_4 & {40{sel[4]}});
    result = result | (input_5 & {40{sel[5]}});
    MUX1HOT_v_40_6_2 = result;
  end
  endfunction


  function automatic [39:0] MUX1HOT_v_40_7_2;
    input [39:0] input_6;
    input [39:0] input_5;
    input [39:0] input_4;
    input [39:0] input_3;
    input [39:0] input_2;
    input [39:0] input_1;
    input [39:0] input_0;
    input [6:0] sel;
    reg [39:0] result;
  begin
    result = input_0 & {40{sel[0]}};
    result = result | (input_1 & {40{sel[1]}});
    result = result | (input_2 & {40{sel[2]}});
    result = result | (input_3 & {40{sel[3]}});
    result = result | (input_4 & {40{sel[4]}});
    result = result | (input_5 & {40{sel[5]}});
    result = result | (input_6 & {40{sel[6]}});
    MUX1HOT_v_40_7_2 = result;
  end
  endfunction


  function automatic [39:0] MUX1HOT_v_40_8_2;
    input [39:0] input_7;
    input [39:0] input_6;
    input [39:0] input_5;
    input [39:0] input_4;
    input [39:0] input_3;
    input [39:0] input_2;
    input [39:0] input_1;
    input [39:0] input_0;
    input [7:0] sel;
    reg [39:0] result;
  begin
    result = input_0 & {40{sel[0]}};
    result = result | (input_1 & {40{sel[1]}});
    result = result | (input_2 & {40{sel[2]}});
    result = result | (input_3 & {40{sel[3]}});
    result = result | (input_4 & {40{sel[4]}});
    result = result | (input_5 & {40{sel[5]}});
    result = result | (input_6 & {40{sel[6]}});
    result = result | (input_7 & {40{sel[7]}});
    MUX1HOT_v_40_8_2 = result;
  end
  endfunction


  function automatic [39:0] MUX1HOT_v_40_9_2;
    input [39:0] input_8;
    input [39:0] input_7;
    input [39:0] input_6;
    input [39:0] input_5;
    input [39:0] input_4;
    input [39:0] input_3;
    input [39:0] input_2;
    input [39:0] input_1;
    input [39:0] input_0;
    input [8:0] sel;
    reg [39:0] result;
  begin
    result = input_0 & {40{sel[0]}};
    result = result | (input_1 & {40{sel[1]}});
    result = result | (input_2 & {40{sel[2]}});
    result = result | (input_3 & {40{sel[3]}});
    result = result | (input_4 & {40{sel[4]}});
    result = result | (input_5 & {40{sel[5]}});
    result = result | (input_6 & {40{sel[6]}});
    result = result | (input_7 & {40{sel[7]}});
    result = result | (input_8 & {40{sel[8]}});
    MUX1HOT_v_40_9_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_5_2;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [4:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    MUX1HOT_v_4_5_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_6_2;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [5:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    MUX1HOT_v_4_6_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_6_2;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [5:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    MUX1HOT_v_5_6_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_7_2;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [6:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    MUX1HOT_v_5_7_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_6_2;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [5:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    MUX1HOT_v_6_6_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_7_2;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [6:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    result = result | (input_4 & {7{sel[4]}});
    result = result | (input_5 & {7{sel[5]}});
    result = result | (input_6 & {7{sel[6]}});
    MUX1HOT_v_7_7_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_4_2;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [3:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    MUX1HOT_v_8_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_6_2;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [5:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    MUX1HOT_v_8_6_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_7_2;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [6:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    MUX1HOT_v_8_7_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_8_2;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [7:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    result = result | (input_7 & {8{sel[7]}});
    MUX1HOT_v_8_8_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_9_2;
    input [7:0] input_8;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [8:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    result = result | (input_7 & {8{sel[7]}});
    result = result | (input_8 & {8{sel[8]}});
    MUX1HOT_v_8_9_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_16_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input  input_4;
    input  input_5;
    input  input_6;
    input  input_7;
    input  input_8;
    input  input_9;
    input  input_10;
    input  input_11;
    input  input_12;
    input  input_13;
    input  input_14;
    input  input_15;
    input [3:0] sel;
    reg  result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_s_1_16_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_4_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input [1:0] sel;
    reg  result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_8_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input  input_4;
    input  input_5;
    input  input_6;
    input  input_7;
    input [2:0] sel;
    reg  result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_s_1_8_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_16_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [11:0] input_2;
    input [11:0] input_3;
    input [11:0] input_4;
    input [11:0] input_5;
    input [11:0] input_6;
    input [11:0] input_7;
    input [11:0] input_8;
    input [11:0] input_9;
    input [11:0] input_10;
    input [11:0] input_11;
    input [11:0] input_12;
    input [11:0] input_13;
    input [11:0] input_14;
    input [11:0] input_15;
    input [3:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_12_16_2 = result;
  end
  endfunction


  function automatic [12:0] MUX_v_13_2_2;
    input [12:0] input_0;
    input [12:0] input_1;
    input  sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_16_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [13:0] input_2;
    input [13:0] input_3;
    input [13:0] input_4;
    input [13:0] input_5;
    input [13:0] input_6;
    input [13:0] input_7;
    input [13:0] input_8;
    input [13:0] input_9;
    input [13:0] input_10;
    input [13:0] input_11;
    input [13:0] input_12;
    input [13:0] input_13;
    input [13:0] input_14;
    input [13:0] input_15;
    input [3:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_14_16_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input  sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_16_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [3:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_16_16_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [22:0] MUX_v_23_16_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [22:0] input_2;
    input [22:0] input_3;
    input [22:0] input_4;
    input [22:0] input_5;
    input [22:0] input_6;
    input [22:0] input_7;
    input [22:0] input_8;
    input [22:0] input_9;
    input [22:0] input_10;
    input [22:0] input_11;
    input [22:0] input_12;
    input [22:0] input_13;
    input [22:0] input_14;
    input [22:0] input_15;
    input [3:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_23_16_2 = result;
  end
  endfunction


  function automatic [23:0] MUX_v_24_16_2;
    input [23:0] input_0;
    input [23:0] input_1;
    input [23:0] input_2;
    input [23:0] input_3;
    input [23:0] input_4;
    input [23:0] input_5;
    input [23:0] input_6;
    input [23:0] input_7;
    input [23:0] input_8;
    input [23:0] input_9;
    input [23:0] input_10;
    input [23:0] input_11;
    input [23:0] input_12;
    input [23:0] input_13;
    input [23:0] input_14;
    input [23:0] input_15;
    input [3:0] sel;
    reg [23:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_24_16_2 = result;
  end
  endfunction


  function automatic [23:0] MUX_v_24_2_2;
    input [23:0] input_0;
    input [23:0] input_1;
    input  sel;
    reg [23:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_24_2_2 = result;
  end
  endfunction


  function automatic [23:0] MUX_v_24_8_2;
    input [23:0] input_0;
    input [23:0] input_1;
    input [23:0] input_2;
    input [23:0] input_3;
    input [23:0] input_4;
    input [23:0] input_5;
    input [23:0] input_6;
    input [23:0] input_7;
    input [2:0] sel;
    reg [23:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_24_8_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_4_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [1:0] input_2;
    input [1:0] input_3;
    input [1:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_2_4_2 = result;
  end
  endfunction


  function automatic [33:0] MUX_v_34_2_2;
    input [33:0] input_0;
    input [33:0] input_1;
    input  sel;
    reg [33:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_34_2_2 = result;
  end
  endfunction


  function automatic [34:0] MUX_v_35_2_2;
    input [34:0] input_0;
    input [34:0] input_1;
    input  sel;
    reg [34:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_35_2_2 = result;
  end
  endfunction


  function automatic [38:0] MUX_v_39_16_2;
    input [38:0] input_0;
    input [38:0] input_1;
    input [38:0] input_2;
    input [38:0] input_3;
    input [38:0] input_4;
    input [38:0] input_5;
    input [38:0] input_6;
    input [38:0] input_7;
    input [38:0] input_8;
    input [38:0] input_9;
    input [38:0] input_10;
    input [38:0] input_11;
    input [38:0] input_12;
    input [38:0] input_13;
    input [38:0] input_14;
    input [38:0] input_15;
    input [3:0] sel;
    reg [38:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_39_16_2 = result;
  end
  endfunction


  function automatic [38:0] MUX_v_39_2_2;
    input [38:0] input_0;
    input [38:0] input_1;
    input  sel;
    reg [38:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_39_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_16_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [2:0] input_4;
    input [2:0] input_5;
    input [2:0] input_6;
    input [2:0] input_7;
    input [2:0] input_8;
    input [2:0] input_9;
    input [2:0] input_10;
    input [2:0] input_11;
    input [2:0] input_12;
    input [2:0] input_13;
    input [2:0] input_14;
    input [2:0] input_15;
    input [3:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_3_16_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_8_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [2:0] input_4;
    input [2:0] input_5;
    input [2:0] input_6;
    input [2:0] input_7;
    input [2:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_3_8_2 = result;
  end
  endfunction


  function automatic [39:0] MUX_v_40_12_2;
    input [39:0] input_0;
    input [39:0] input_1;
    input [39:0] input_2;
    input [39:0] input_3;
    input [39:0] input_4;
    input [39:0] input_5;
    input [39:0] input_6;
    input [39:0] input_7;
    input [39:0] input_8;
    input [39:0] input_9;
    input [39:0] input_10;
    input [39:0] input_11;
    input [3:0] sel;
    reg [39:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      default : begin
        result = input_11;
      end
    endcase
    MUX_v_40_12_2 = result;
  end
  endfunction


  function automatic [39:0] MUX_v_40_15_2;
    input [39:0] input_0;
    input [39:0] input_1;
    input [39:0] input_2;
    input [39:0] input_3;
    input [39:0] input_4;
    input [39:0] input_5;
    input [39:0] input_6;
    input [39:0] input_7;
    input [39:0] input_8;
    input [39:0] input_9;
    input [39:0] input_10;
    input [39:0] input_11;
    input [39:0] input_12;
    input [39:0] input_13;
    input [39:0] input_14;
    input [3:0] sel;
    reg [39:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      default : begin
        result = input_14;
      end
    endcase
    MUX_v_40_15_2 = result;
  end
  endfunction


  function automatic [39:0] MUX_v_40_16_2;
    input [39:0] input_0;
    input [39:0] input_1;
    input [39:0] input_2;
    input [39:0] input_3;
    input [39:0] input_4;
    input [39:0] input_5;
    input [39:0] input_6;
    input [39:0] input_7;
    input [39:0] input_8;
    input [39:0] input_9;
    input [39:0] input_10;
    input [39:0] input_11;
    input [39:0] input_12;
    input [39:0] input_13;
    input [39:0] input_14;
    input [39:0] input_15;
    input [3:0] sel;
    reg [39:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_40_16_2 = result;
  end
  endfunction


  function automatic [39:0] MUX_v_40_2_2;
    input [39:0] input_0;
    input [39:0] input_1;
    input  sel;
    reg [39:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_40_2_2 = result;
  end
  endfunction


  function automatic [39:0] MUX_v_40_4_2;
    input [39:0] input_0;
    input [39:0] input_1;
    input [39:0] input_2;
    input [39:0] input_3;
    input [1:0] sel;
    reg [39:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_40_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [52:0] MUX_v_53_2_2;
    input [52:0] input_0;
    input [52:0] input_1;
    input  sel;
    reg [52:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_53_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_16_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [7:0] input_10;
    input [7:0] input_11;
    input [7:0] input_12;
    input [7:0] input_13;
    input [7:0] input_14;
    input [7:0] input_15;
    input [3:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_8_16_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_8_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_16_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [8:0] input_2;
    input [8:0] input_3;
    input [8:0] input_4;
    input [8:0] input_5;
    input [8:0] input_6;
    input [8:0] input_7;
    input [8:0] input_8;
    input [8:0] input_9;
    input [8:0] input_10;
    input [8:0] input_11;
    input [8:0] input_12;
    input [8:0] input_13;
    input [8:0] input_14;
    input [8:0] input_15;
    input [3:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_9_16_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_26_1_25;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 25;
    readslicef_26_1_25 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_3_1_2;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_3_1_2 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_41_1_40;
    input [40:0] vector;
    reg [40:0] tmp;
  begin
    tmp = vector >> 40;
    readslicef_41_1_40 = tmp[0:0];
  end
  endfunction


  function automatic [39:0] readslicef_41_40_1;
    input [40:0] vector;
    reg [40:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_41_40_1 = tmp[39:0];
  end
  endfunction


  function automatic [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function automatic [39:0] readslicef_56_40_16;
    input [55:0] vector;
    reg [55:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_56_40_16 = tmp[39:0];
  end
  endfunction


  function automatic [43:0] readslicef_72_44_28;
    input [71:0] vector;
    reg [71:0] tmp;
  begin
    tmp = vector >> 28;
    readslicef_72_44_28 = tmp[43:0];
  end
  endfunction


  function automatic [14:0] signext_15_1;
    input  vector;
  begin
    signext_15_1= {{14{vector}}, vector};
  end
  endfunction


  function automatic [15:0] signext_16_14;
    input [13:0] vector;
  begin
    signext_16_14= {{2{vector[13]}}, vector};
  end
  endfunction


  function automatic [21:0] signext_22_1;
    input  vector;
  begin
    signext_22_1= {{21{vector}}, vector};
  end
  endfunction


  function automatic [23:0] signext_24_4;
    input [3:0] vector;
  begin
    signext_24_4= {{20{vector[3]}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input  vector;
  begin
    signext_2_1= {{1{vector}}, vector};
  end
  endfunction


  function automatic [38:0] signext_39_33;
    input [32:0] vector;
  begin
    signext_39_33= {{6{vector[32]}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_1;
    input  vector;
  begin
    signext_3_1= {{2{vector}}, vector};
  end
  endfunction


  function automatic [39:0] signext_40_30;
    input [29:0] vector;
  begin
    signext_40_30= {{10{vector[29]}}, vector};
  end
  endfunction


  function automatic [52:0] signext_53_52;
    input [51:0] vector;
  begin
    signext_53_52= {{1{vector[51]}}, vector};
  end
  endfunction


  function automatic [5:0] signext_6_1;
    input  vector;
  begin
    signext_6_1= {{5{vector}}, vector};
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input  vector;
  begin
    signext_7_1= {{6{vector}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_8_24 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_24 = {{16{vector[7]}}, vector};
  end
  endfunction


  function automatic [40:0] conv_s2s_40_41 ;
    input [39:0]  vector ;
  begin
    conv_s2s_40_41 = {vector[39], vector};
  end
  endfunction


  function automatic [40:0] conv_s2u_40_41 ;
    input [39:0]  vector ;
  begin
    conv_s2u_40_41 = {vector[39], vector};
  end
  endfunction


  function automatic [35:0] conv_u2s_1_36 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_36 = {{35{1'b0}}, vector};
  end
  endfunction


  function automatic [38:0] conv_u2s_1_39 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_39 = {{38{1'b0}}, vector};
  end
  endfunction


  function automatic [2:0] conv_u2s_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2s_2_3 =  {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [16:0] conv_u2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2s_16_17 =  {1'b0, vector};
  end
  endfunction


  function automatic [20:0] conv_u2s_20_21 ;
    input [19:0]  vector ;
  begin
    conv_u2s_20_21 =  {1'b0, vector};
  end
  endfunction


  function automatic [35:0] conv_u2s_35_36 ;
    input [34:0]  vector ;
  begin
    conv_u2s_35_36 =  {1'b0, vector};
  end
  endfunction


  function automatic [39:0] conv_u2s_39_40 ;
    input [38:0]  vector ;
  begin
    conv_u2s_39_40 =  {1'b0, vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_3 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    dut
// ------------------------------------------------------------------


module dut (
  clk, en, rst, strm_in_rsc_dat, strm_in_rsc_vld, strm_in_rsc_rdy, strm_out_rsc_dat,
      strm_out_rsc_vld, strm_out_rsc_rdy
);
  input clk;
  input en;
  input rst;
  input [31:0] strm_in_rsc_dat;
  input strm_in_rsc_vld;
  output strm_in_rsc_rdy;
  output [31:0] strm_out_rsc_dat;
  output strm_out_rsc_vld;
  input strm_out_rsc_rdy;


  // Interconnect Declarations
  wire attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d;
  wire [39:0] attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d;
  wire [39:0] attention_2_1_16_16_4_4_k_cache_upd_rsci_q_d;
  wire [5:0] attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d;
  wire [5:0] attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d;
  wire [39:0] attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d;
  wire [39:0] attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d;
  wire [5:0] attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d;
  wire [5:0] attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d;
  wire [39:0] attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d;
  wire [5:0] attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d;
  wire [5:0] attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d;
  wire [71:0] rms_norm_16_div_cmp_a;
  wire [60:0] rms_norm_16_div_cmp_b;
  wire [71:0] rms_norm_16_div_cmp_z;
  wire attention_2_1_16_16_4_4_k_cache_upd_rsc_clken;
  wire [39:0] attention_2_1_16_16_4_4_k_cache_upd_rsc_q;
  wire attention_2_1_16_16_4_4_k_cache_upd_rsc_re;
  wire [5:0] attention_2_1_16_16_4_4_k_cache_upd_rsc_radr;
  wire attention_2_1_16_16_4_4_k_cache_upd_rsc_we;
  wire [39:0] attention_2_1_16_16_4_4_k_cache_upd_rsc_d;
  wire [5:0] attention_2_1_16_16_4_4_k_cache_upd_rsc_wadr;
  wire attention_2_1_16_16_4_4_v_cache_upd_rsc_clken;
  wire [39:0] attention_2_1_16_16_4_4_v_cache_upd_rsc_q;
  wire attention_2_1_16_16_4_4_v_cache_upd_rsc_re;
  wire [5:0] attention_2_1_16_16_4_4_v_cache_upd_rsc_radr;
  wire attention_2_1_16_16_4_4_v_cache_upd_rsc_we;
  wire [39:0] attention_2_1_16_16_4_4_v_cache_upd_rsc_d;
  wire [5:0] attention_2_1_16_16_4_4_v_cache_upd_rsc_wadr;
  wire attention_2_1_16_16_4_4_k_proj_transposed_rsc_clken;
  wire [39:0] attention_2_1_16_16_4_4_k_proj_transposed_rsc_q;
  wire attention_2_1_16_16_4_4_k_proj_transposed_rsc_re;
  wire [5:0] attention_2_1_16_16_4_4_k_proj_transposed_rsc_radr;
  wire attention_2_1_16_16_4_4_k_proj_transposed_rsc_we;
  wire [39:0] attention_2_1_16_16_4_4_k_proj_transposed_rsc_d;
  wire [5:0] attention_2_1_16_16_4_4_k_proj_transposed_rsc_wadr;
  wire attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_iff;
  wire attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_iff;
  wire attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_iff;
  wire attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_iff;
  wire attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  mgc_div #(.width_a(32'sd72),
  .width_b(32'sd61),
  .signd(32'sd1)) rms_norm_16_div_cmp (
      .a(rms_norm_16_div_cmp_a),
      .b(rms_norm_16_div_cmp_b),
      .z(rms_norm_16_div_cmp_z)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd6),
  .data_width(32'sd40),
  .depth(32'sd48),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) attention_2_1_16_16_4_4_k_cache_upd_rsc_comp
      (
      .clk(clk),
      .clken(attention_2_1_16_16_4_4_k_cache_upd_rsc_clken),
      .d(attention_2_1_16_16_4_4_k_cache_upd_rsc_d),
      .q(attention_2_1_16_16_4_4_k_cache_upd_rsc_q),
      .radr(attention_2_1_16_16_4_4_k_cache_upd_rsc_radr),
      .re(attention_2_1_16_16_4_4_k_cache_upd_rsc_re),
      .wadr(attention_2_1_16_16_4_4_k_cache_upd_rsc_wadr),
      .we(attention_2_1_16_16_4_4_k_cache_upd_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd6),
  .data_width(32'sd40),
  .depth(32'sd48),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) attention_2_1_16_16_4_4_v_cache_upd_rsc_comp
      (
      .clk(clk),
      .clken(attention_2_1_16_16_4_4_v_cache_upd_rsc_clken),
      .d(attention_2_1_16_16_4_4_v_cache_upd_rsc_d),
      .q(attention_2_1_16_16_4_4_v_cache_upd_rsc_q),
      .radr(attention_2_1_16_16_4_4_v_cache_upd_rsc_radr),
      .re(attention_2_1_16_16_4_4_v_cache_upd_rsc_re),
      .wadr(attention_2_1_16_16_4_4_v_cache_upd_rsc_wadr),
      .we(attention_2_1_16_16_4_4_v_cache_upd_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd6),
  .data_width(32'sd40),
  .depth(32'sd48),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) attention_2_1_16_16_4_4_k_proj_transposed_rsc_comp
      (
      .clk(clk),
      .clken(attention_2_1_16_16_4_4_k_proj_transposed_rsc_clken),
      .d(attention_2_1_16_16_4_4_k_proj_transposed_rsc_d),
      .q(attention_2_1_16_16_4_4_k_proj_transposed_rsc_q),
      .radr(attention_2_1_16_16_4_4_k_proj_transposed_rsc_radr),
      .re(attention_2_1_16_16_4_4_k_proj_transposed_rsc_re),
      .wadr(attention_2_1_16_16_4_4_k_proj_transposed_rsc_wadr),
      .we(attention_2_1_16_16_4_4_k_proj_transposed_rsc_we)
    );
  dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_14_6_40_48_1_48_40_1_gen attention_2_1_16_16_4_4_k_cache_upd_rsci
      (
      .clken(attention_2_1_16_16_4_4_k_cache_upd_rsc_clken),
      .q(attention_2_1_16_16_4_4_k_cache_upd_rsc_q),
      .re(attention_2_1_16_16_4_4_k_cache_upd_rsc_re),
      .radr(attention_2_1_16_16_4_4_k_cache_upd_rsc_radr),
      .we(attention_2_1_16_16_4_4_k_cache_upd_rsc_we),
      .d(attention_2_1_16_16_4_4_k_cache_upd_rsc_d),
      .wadr(attention_2_1_16_16_4_4_k_cache_upd_rsc_wadr),
      .clken_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d),
      .d_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d),
      .q_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_q_d),
      .radr_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d),
      .re_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_iff),
      .wadr_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d),
      .we_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_iff)
    );
  dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_15_6_40_48_1_48_40_1_gen attention_2_1_16_16_4_4_v_cache_upd_rsci
      (
      .clken(attention_2_1_16_16_4_4_v_cache_upd_rsc_clken),
      .q(attention_2_1_16_16_4_4_v_cache_upd_rsc_q),
      .re(attention_2_1_16_16_4_4_v_cache_upd_rsc_re),
      .radr(attention_2_1_16_16_4_4_v_cache_upd_rsc_radr),
      .we(attention_2_1_16_16_4_4_v_cache_upd_rsc_we),
      .d(attention_2_1_16_16_4_4_v_cache_upd_rsc_d),
      .wadr(attention_2_1_16_16_4_4_v_cache_upd_rsc_wadr),
      .clken_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d),
      .d_d(attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d),
      .q_d(attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d),
      .radr_d(attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d),
      .re_d(attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_iff),
      .wadr_d(attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d),
      .we_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_iff)
    );
  dut_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_16_6_40_48_1_48_40_1_gen attention_2_1_16_16_4_4_k_proj_transposed_rsci
      (
      .clken(attention_2_1_16_16_4_4_k_proj_transposed_rsc_clken),
      .q(attention_2_1_16_16_4_4_k_proj_transposed_rsc_q),
      .re(attention_2_1_16_16_4_4_k_proj_transposed_rsc_re),
      .radr(attention_2_1_16_16_4_4_k_proj_transposed_rsc_radr),
      .we(attention_2_1_16_16_4_4_k_proj_transposed_rsc_we),
      .d(attention_2_1_16_16_4_4_k_proj_transposed_rsc_d),
      .wadr(attention_2_1_16_16_4_4_k_proj_transposed_rsc_wadr),
      .clken_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d),
      .d_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_q_d),
      .q_d(attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d),
      .radr_d(attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d),
      .re_d(attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_iff),
      .wadr_d(attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d),
      .we_d(attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_iff)
    );
  dut_core dut_core_inst (
      .clk(clk),
      .en(en),
      .rst(rst),
      .strm_in_rsc_dat(strm_in_rsc_dat),
      .strm_in_rsc_vld(strm_in_rsc_vld),
      .strm_in_rsc_rdy(strm_in_rsc_rdy),
      .strm_out_rsc_dat(strm_out_rsc_dat),
      .strm_out_rsc_vld(strm_out_rsc_vld),
      .strm_out_rsc_rdy(strm_out_rsc_rdy),
      .attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_clken_d),
      .attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_d_d),
      .attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_radr_d),
      .attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d(attention_2_1_16_16_4_4_k_cache_upd_rsci_wadr_d),
      .attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d(attention_2_1_16_16_4_4_v_cache_upd_rsci_d_d),
      .attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d(attention_2_1_16_16_4_4_v_cache_upd_rsci_q_d),
      .attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d(attention_2_1_16_16_4_4_v_cache_upd_rsci_radr_d),
      .attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d(attention_2_1_16_16_4_4_v_cache_upd_rsci_wadr_d),
      .attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d(attention_2_1_16_16_4_4_k_proj_transposed_rsci_q_d),
      .attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d(attention_2_1_16_16_4_4_k_proj_transposed_rsci_radr_d),
      .attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d(attention_2_1_16_16_4_4_k_proj_transposed_rsci_wadr_d),
      .rms_norm_16_div_cmp_a(rms_norm_16_div_cmp_a),
      .rms_norm_16_div_cmp_b(rms_norm_16_div_cmp_b),
      .rms_norm_16_div_cmp_z(rms_norm_16_div_cmp_z),
      .attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_pff(attention_2_1_16_16_4_4_k_cache_upd_rsci_re_d_iff),
      .attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_pff(attention_2_1_16_16_4_4_k_cache_upd_rsci_we_d_iff),
      .attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_pff(attention_2_1_16_16_4_4_v_cache_upd_rsci_re_d_iff),
      .attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_pff(attention_2_1_16_16_4_4_k_proj_transposed_rsci_re_d_iff),
      .attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_pff(attention_2_1_16_16_4_4_k_proj_transposed_rsci_we_d_iff)
    );
endmodule



